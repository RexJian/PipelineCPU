//Precision RTL Synthesis 64-bit 2023.1.0.14 (Production Release) Fri Feb 17 02:47:53 PST 2023
//
//           This material contains trade secrets or otherwise confidential
//           information owned by Siemens Industry Software Inc. or its    
//           affiliates (collectively, "Siemens"), or its licensors. Access to
//           and use of this information is strictly limited as set forth    
//           in the Customer's applicable agreements with Siemens.           
//
//                            Unpublished work. Copyright 2023 Siemens               
//
//Running on Linux runner@043ec5d9170f #201-Ubuntu SMP Thu Mar 28 15:39:01 UTC 2024 5.4.0-181-generic x86_64
//
//
// Verilog description for cell main, 
//

module main ( CLK, EN, CLR_N, Addr, Alu_D1, Y, Ex_Alu_R, Write_D, stall, 
              condition_met, Rs, Rt, Rd ) ;

    input CLK ;
    input EN ;
    input CLR_N ;
    output [31:0]Addr ;
    output [31:0]Alu_D1 ;
    output [31:0]Y ;
    output [31:0]Ex_Alu_R ;
    output [31:0]Write_D ;
    output stall ;
    output condition_met ;
    output [4:0]Rs ;
    output [4:0]Rt ;
    output [4:0]Rd ;

    wire [31:0]Addr_1_0;
    wire \Rs_1_0(2)  , \Rs_1_0(1)  , \Rs_1_0(0)  , \Rt_1_0(2)  , \Rt_1_0(1)  , 
         \Rt_1_0(0)  , \Rd_1_0(2)  , \Rd_1_0(1)  , \Rd_1_0(0)  ;
    wire \Pc_Add4(31)  , \Pc_Add4(30)  , \Pc_Add4(29)  , \Pc_Add4(28)  , 
         \Pc_Add4(27)  , \Pc_Add4(26)  , \Pc_Add4(25)  , \Pc_Add4(24)  , 
         \Pc_Add4(23)  , \Pc_Add4(22)  , \Pc_Add4(21)  , \Pc_Add4(20)  , 
         \Pc_Add4(19)  , \Pc_Add4(18)  , \Pc_Add4(17)  , \Pc_Add4(16)  , 
         \Pc_Add4(15)  , \Pc_Add4(14)  , \Pc_Add4(13)  , \Pc_Add4(12)  , 
         \Pc_Add4(11)  , \Pc_Add4(10)  , \Pc_Add4(9)  , \Pc_Add4(8)  , 
         \Pc_Add4(7)  , \Pc_Add4(6)  , \Pc_Add4(5)  , \Pc_Add4(4)  , 
         \Pc_Add4(3)  , \Pc_Add4(2)  ;
    wire [31:0]Id_Pc_Add4;
    wire \Id_Inst(29)  , \Id_Inst(28)  , \Id_Inst(26)  , \Id_Extimm(13)  , 
         \Id_Extimm(12)  , \Id_Extimm(11)  , \Id_Extimm(4)  ;
    wire \Id_Extimm(3)  , \Id_Extimm(2)  , \Id_Extimm(1)  , \Id_Extimm(0)  ;
    wire [31:0]Ex_D1;
    wire [31:0]Ex_D2;
    wire \Ex_Extimm(13)  , \Ex_Extimm(0)  ;
    wire [31:0]Mem_Alu_R;
    wire [31:0]Mem_D2;
    wire [31:0]Wb_D;
    wire [31:0]Wb_Alu_R;
    wire \Instruction(31)  , \Instruction(29)  , \Instruction(28)  , 
         \Instruction(23)  , \Instruction(22)  , \Instruction(21)  , 
         \Instruction(18)  , \Instruction(17)  , \Instruction(16)  , 
         \Instruction(13)  , \Instruction(12)  , \Instruction(11)  , 
         \Instruction(4)  , \Instruction(3)  , \Instruction(2)  , 
         \Instruction(1)  , \Instruction(0)  ;
    wire [31:0]Next_Addr;
    wire \Ex_Op(0)  ;
    wire [2:0]Ex_Rd;
    wire [2:0]Mem_Rd;
    wire Ex_Z;
    wire Ex_Wreg, Ex_Reg2reg, Ex_Wmem, Ex_Aluqb, Mem_Wreg, Mem_Reg2reg, Wb_Wreg, 
         Wb_Reg2reg;
    wire [1:0]Ex_Fwd_A;
    wire [1:0]Ex_Fwd_B;
    wire [2:0]Ex_Aluc;
    wire Mem_Wmem, nx759z33, nx759z31, nx759z30, nx759z29, nx759z28, nx759z27, 
         nx759z26, nx759z25, nx759z24, nx759z23, nx759z22, nx759z21, nx759z20, 
         nx759z19, nx759z18, nx759z17, nx759z16, nx759z15, nx759z14, nx759z13, 
         nx759z12, nx759z11, nx759z10, nx759z9, nx759z8, nx759z7, nx759z6, 
         nx759z5, nx759z4, nx759z3, nx759z2, nx759z1, nx759z66, nx759z64, 
         nx759z63, nx759z62, nx759z61, nx759z60, nx759z59, nx759z58, nx759z57, 
         nx759z56, nx759z55, nx759z54, nx759z53, nx759z52, nx759z51, nx759z50, 
         nx759z49, nx759z48, nx759z47, nx759z46, nx759z45, nx759z44, nx759z43, 
         nx759z42, nx759z41, nx759z40, nx759z39, nx759z38, nx759z37, nx759z36, 
         nx759z35, nx759z34, nx22656z32, nx22656z31, nx22656z30, nx22656z29, 
         nx22656z28, nx22656z27, nx22656z26, nx22656z25, nx22656z24, nx22656z23, 
         nx22656z22, nx22656z21, nx22656z20, nx22656z19, nx22656z18, nx22656z17, 
         nx22656z16, nx22656z15, nx22656z14, nx22656z13, nx22656z12, nx22656z11, 
         nx22656z10, nx22656z9, nx22656z8, nx22656z7, nx22656z6, nx22656z5, 
         nx22656z4, nx22656z3, nx22656z2, nx22656z1;
    wire CLK_int;
    wire EN_int, CLR_N_int, pc_not_clr_n, nx15902z32, nx57674z45, nx15902z1, 
         nx15902z2, nx15902z3, nx15902z4, nx15902z5, nx15902z6, nx15902z7, 
         nx15902z8, nx15902z9, nx15902z10, nx15902z11, nx15902z12, nx15902z13, 
         nx15902z14, nx15902z15, nx15902z16, nx15902z17, nx15902z18, nx15902z19, 
         nx15902z20, nx15902z21, nx15902z22, nx15902z23, nx15902z24, nx15902z25, 
         nx15902z26, nx15902z27, nx15902z28, nx15902z29, nx15902z30, nx15902z31, 
         nx15902z33, nx10566z1, nx11563z1, nx13559z1, nx14556z1, nx15553z1, 
         nx16550z1, nx17547z1, nx18544z1, nx19541z1, nx20538z1, nx21535z1, 
         nx22532z1, nx24528z1, nx25525z1, nx26522z1, nx27519z1, nx28516z1, 
         nx29513z1, nx30510z1, nx31507z1, nx32504z1, nx33501z1, nx13165z1, 
         nx14162z1, nx15159z1, nx16156z1, nx17153z1, nx18150z1, nx19147z1, 
         nx20144z1, nx21141z1, nx22138z1, nx32823z1, nx33820z1, nx34817z1, 
         nx9585z1, nx10582z1, nx11579z1, nx12576z1, nx13573z1, nx14570z1, 
         nx54097z77, nx54097z76, nx54097z75, nx54097z74, nx54097z73, nx54097z72, 
         nx54097z71, nx54097z70, nx54097z69, nx54097z68, nx54097z67, nx54097z66, 
         nx54097z65, nx54097z64, nx54097z63, nx54097z62, nx54097z61, nx54097z60, 
         nx54097z59, nx54097z58, nx54097z57, nx54097z56, nx54097z55, nx54097z54, 
         nx54097z53, nx54097z52, nx54097z51, nx26565z1, nx27562z1, nx28559z1, 
         nx29556z1, nx30553z1, nx53980z1, nx54977z1, nx55974z1, nx56971z1, 
         nx57968z1, nx58965z1, nx59962z1, nx60959z1, nx61956z1, nx62953z1, 
         nx30993z1, nx31990z1, nx32987z1, nx33984z1, nx34981z1, nx35978z1, 
         nx36975z1, nx37972z1, nx38969z1, nx39966z1, nx41962z1, nx42959z1, 
         nx43956z1, nx44953z1, nx45950z1, nx46947z1, nx47944z1, nx48941z1, 
         nx49938z1, nx50935z1, nx52931z1, nx53928z1, nx3137z1, nx2140z1, 
         nx1143z1, nx146z1, nx64685z1, nx63688z1, nx62691z1, nx61694z1, 
         nx60697z1, nx59700z1, nx29408z1, nx28411z1, nx27414z1, nx26417z1, 
         nx25420z1, nx24423z1, nx23426z1, nx22429z1, nx21432z1, nx20435z1, 
         nx18439z1, nx17442z1, nx16445z1, nx15448z1, nx14451z1, nx13454z1, 
         nx12457z1, nx11460z1, nx10463z1, nx9466z1, nx7470z1, nx6473z1, 
         nx17673z32, nx17673z31, nx17673z30, nx17673z29, nx17673z28, nx17673z27, 
         nx17673z26, nx17673z25, nx17673z24, nx17673z23, nx17673z22, nx17673z21, 
         nx17673z20, nx17673z19, nx17673z18, nx17673z17, nx17673z16, nx17673z15, 
         nx17673z14, nx17673z13, nx17673z12, nx17673z11, nx17673z10, nx17673z9, 
         nx17673z8, nx17673z7, nx17673z6, nx17673z5, nx17673z4, nx17673z3, 
         nx17673z2, nx17673z1, nx57674z37, nx57674z38, nx57674z39, nx57674z40, 
         nx57674z41, nx57674z42, nx57674z43, nx57674z44, nx23941z17, nx54097z29, 
         nx23941z18, nx54097z28, nx57674z30, nx54097z30, nx57674z27, nx54097z31, 
         nx57674z26, nx54097z33, nx57674z25, nx54097z34, nx57674z24, nx54097z35, 
         nx57674z23, nx54097z36, nx57674z22, nx54097z42, nx57674z21, nx54097z48, 
         nx57674z20, nx21854z1, nx57674z19, nx54097z49, nx57674z18, nx54097z45, 
         nx57674z17, nx54097z46, nx57674z16, nx54097z43, nx57674z15, nx54097z50, 
         nx57674z14, nx54097z39, nx57674z13, nx54097z32, nx57674z12, nx54097z47, 
         nx57674z11, nx54097z44, nx57674z10, nx23941z16, nx57674z9, nx57674z36, 
         nx23941z15, nx57674z8, nx57674z35, nx23941z14, nx57674z7, nx54097z40, 
         nx57674z6, nx54097z41, nx57674z5, nx54097z37, nx57674z4, nx54097z38, 
         nx57674z3, nx57674z31, nx23941z7, nx57674z1, nx57674z2, nx23941z1, 
         nx23941z2, nx54097z1, nx63922z1, nx64919z1, nx380z1, nx1377z1, nx2374z1, 
         nx3371z1, nx4368z1, nx5365z1, nx6362z1, nx7359z1, nx47231z1, nx48228z1, 
         nx49225z1, nx50222z1, nx51219z1, nx52216z1, nx53213z1, nx54210z1, 
         nx55207z1, nx56204z1, nx58200z1, nx59197z1, nx60194z1, nx61191z1, 
         nx62188z1, nx63185z1, nx64182z1, nx65179z1, nx640z1, nx1637z1, nx3633z1, 
         nx4630z1, nx57674z32, nx23941z8, nx23941z3, nx57674z33, nx23941z9, 
         nx23941z4, nx57674z34, nx23941z10, nx23941z5, nx23941z6, nx23941z11, 
         nx58593z1, nx57674z28, nx57674z29, nx23941z12, nx759z65, nx59962z2, 
         nx759z32, nx28580z1, nx4583z1, nx42977z1, nx42977z2, nx60794z1, 
         nx17673z33, nx54097z2, nx23941z13, nx54097z3, nx54097z4, nx54097z5, 
         nx54097z6, nx54097z7, nx54097z8, nx54097z9, nx54097z10, nx54097z11, 
         nx54097z12, nx54097z13, nx54097z14, nx54097z15, nx54097z16, nx54097z17, 
         nx54097z18, nx54097z19, nx54097z20, nx54097z21, nx54097z22, nx54097z23, 
         nx54097z24, nx54097z25, nx54097z26, nx54097z27;
    wire [213:0] \$dummy ;




    ram_dq_32_0 register (.wr_data1 ({nx17673z1,nx17673z2,nx17673z3,nx17673z4,
                nx17673z5,nx17673z6,nx17673z7,nx17673z8,nx17673z9,nx17673z10,
                nx17673z11,nx17673z12,nx17673z13,nx17673z14,nx17673z15,
                nx17673z16,nx17673z17,nx17673z18,nx17673z19,nx17673z20,
                nx17673z21,nx17673z22,nx17673z23,nx17673z24,nx17673z25,
                nx17673z26,nx17673z27,nx17673z28,nx17673z29,nx17673z30,
                nx17673z31,nx17673z32}), .addr1 ({\$dummy [0],\$dummy [1],
                \Rd_1_0(2)  ,\Rd_1_0(1)  ,\Rd_1_0(0)  }), .wr_clk1 (CLK_int), .wr_ena1 (
                nx17673z33), .rd_data2 ({nx759z1,nx759z2,nx759z3,nx759z4,nx759z5
                ,nx759z6,nx759z7,nx759z8,nx759z9,nx759z10,nx759z11,nx759z12,
                nx759z13,nx759z14,nx759z15,nx759z16,nx759z17,nx759z18,nx759z19,
                nx759z20,nx759z21,nx759z22,nx759z23,nx759z24,nx759z25,nx759z26,
                nx759z27,nx759z28,nx759z29,nx759z30,nx759z31,nx759z33}), .addr2 (
                {\$dummy [2],\$dummy [3],\Rs_1_0(2)  ,\Rs_1_0(1)  ,\Rs_1_0(0)  }
                ), .rd_data3 ({nx759z34,nx759z35,nx759z36,nx759z37,nx759z38,
                nx759z39,nx759z40,nx759z41,nx759z42,nx759z43,nx759z44,nx759z45,
                nx759z46,nx759z47,nx759z48,nx759z49,nx759z50,nx759z51,nx759z52,
                nx759z53,nx759z54,nx759z55,nx759z56,nx759z57,nx759z58,nx759z59,
                nx759z60,nx759z61,nx759z62,nx759z63,nx759z64,nx759z66}), .addr3 (
                {\$dummy [4],\$dummy [5],\Rt_1_0(2)  ,\Rt_1_0(1)  ,\Rt_1_0(0)  }
                )) ;
    ram_dq_32_1 ROM (.wr_data1 ({Mem_D2[31],Mem_D2[30],Mem_D2[29],Mem_D2[28],
                Mem_D2[27],Mem_D2[26],Mem_D2[25],Mem_D2[24],Mem_D2[23],
                Mem_D2[22],Mem_D2[21],Mem_D2[20],Mem_D2[19],Mem_D2[18],
                Mem_D2[17],Mem_D2[16],Mem_D2[15],Mem_D2[14],Mem_D2[13],
                Mem_D2[12],Mem_D2[11],Mem_D2[10],Mem_D2[9],Mem_D2[8],Mem_D2[7],
                Mem_D2[6],Mem_D2[5],Mem_D2[4],Mem_D2[3],Mem_D2[2],Mem_D2[1],
                Mem_D2[0]}), .addr1 ({Mem_Alu_R[6],Mem_Alu_R[5],Mem_Alu_R[4],
                Mem_Alu_R[3],Mem_Alu_R[2]}), .wr_clk1 (CLK_int), .wr_ena1 (
                nx60794z1), .rd_data2 ({nx22656z1,nx22656z2,nx22656z3,nx22656z4,
                nx22656z5,nx22656z6,nx22656z7,nx22656z8,nx22656z9,nx22656z10,
                nx22656z11,nx22656z12,nx22656z13,nx22656z14,nx22656z15,
                nx22656z16,nx22656z17,nx22656z18,nx22656z19,nx22656z20,
                nx22656z21,nx22656z22,nx22656z23,nx22656z24,nx22656z25,
                nx22656z26,nx22656z27,nx22656z28,nx22656z29,nx22656z30,
                nx22656z31,nx22656z32})) ;
    inc_30_0 pc_add4_PC_Add4_inc30_0 (.a ({Addr_1_0[31],Addr_1_0[30],
             Addr_1_0[29],Addr_1_0[28],Addr_1_0[27],Addr_1_0[26],Addr_1_0[25],
             Addr_1_0[24],Addr_1_0[23],Addr_1_0[22],Addr_1_0[21],Addr_1_0[20],
             Addr_1_0[19],Addr_1_0[18],Addr_1_0[17],Addr_1_0[16],Addr_1_0[15],
             Addr_1_0[14],Addr_1_0[13],Addr_1_0[12],Addr_1_0[11],Addr_1_0[10],
             Addr_1_0[9],Addr_1_0[8],Addr_1_0[7],Addr_1_0[6],Addr_1_0[5],
             Addr_1_0[4],Addr_1_0[3],Addr_1_0[2]}), .d ({\Pc_Add4(31)  ,
             \Pc_Add4(30)  ,\Pc_Add4(29)  ,\Pc_Add4(28)  ,\Pc_Add4(27)  ,
             \Pc_Add4(26)  ,\Pc_Add4(25)  ,\Pc_Add4(24)  ,\Pc_Add4(23)  ,
             \Pc_Add4(22)  ,\Pc_Add4(21)  ,\Pc_Add4(20)  ,\Pc_Add4(19)  ,
             \Pc_Add4(18)  ,\Pc_Add4(17)  ,\Pc_Add4(16)  ,\Pc_Add4(15)  ,
             \Pc_Add4(14)  ,\Pc_Add4(13)  ,\Pc_Add4(12)  ,\Pc_Add4(11)  ,
             \Pc_Add4(10)  ,\Pc_Add4(9)  ,\Pc_Add4(8)  ,\Pc_Add4(7)  ,
             \Pc_Add4(6)  ,\Pc_Add4(5)  ,\Pc_Add4(4)  ,\Pc_Add4(3)  ,
             \Pc_Add4(2)  })) ;
    FDRE \reg_Rs(2)  (.Q (\Rs_1_0(2)  ), .C (CLK_int), .CE (nx42977z1), .D (
         \Instruction(23)  ), .R (nx28580z1)) ;
    FDRE \reg_Rs(1)  (.Q (\Rs_1_0(1)  ), .C (CLK_int), .CE (nx42977z1), .D (
         \Instruction(22)  ), .R (nx28580z1)) ;
    FDRE \reg_Rs(0)  (.Q (\Rs_1_0(0)  ), .C (CLK_int), .CE (nx42977z1), .D (
         \Instruction(21)  ), .R (nx28580z1)) ;
    FDRE \reg_Rt(2)  (.Q (\Rt_1_0(2)  ), .C (CLK_int), .CE (nx42977z1), .D (
         \Instruction(18)  ), .R (nx28580z1)) ;
    FDRE \reg_Rt(1)  (.Q (\Rt_1_0(1)  ), .C (CLK_int), .CE (nx42977z1), .D (
         \Instruction(17)  ), .R (nx28580z1)) ;
    FDRE \reg_Rt(0)  (.Q (\Rt_1_0(0)  ), .C (CLK_int), .CE (nx42977z1), .D (
         \Instruction(16)  ), .R (nx28580z1)) ;
    FDRE \reg_Ex_D1(31)  (.Q (Ex_D1[31]), .C (CLK_int), .CE (EN_int), .D (
         nx6473z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(30)  (.Q (Ex_D1[30]), .C (CLK_int), .CE (EN_int), .D (
         nx7470z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(29)  (.Q (Ex_D1[29]), .C (CLK_int), .CE (EN_int), .D (
         nx9466z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(28)  (.Q (Ex_D1[28]), .C (CLK_int), .CE (EN_int), .D (
         nx10463z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(27)  (.Q (Ex_D1[27]), .C (CLK_int), .CE (EN_int), .D (
         nx11460z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(26)  (.Q (Ex_D1[26]), .C (CLK_int), .CE (EN_int), .D (
         nx12457z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(25)  (.Q (Ex_D1[25]), .C (CLK_int), .CE (EN_int), .D (
         nx13454z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(24)  (.Q (Ex_D1[24]), .C (CLK_int), .CE (EN_int), .D (
         nx14451z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(23)  (.Q (Ex_D1[23]), .C (CLK_int), .CE (EN_int), .D (
         nx15448z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(22)  (.Q (Ex_D1[22]), .C (CLK_int), .CE (EN_int), .D (
         nx16445z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(21)  (.Q (Ex_D1[21]), .C (CLK_int), .CE (EN_int), .D (
         nx17442z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(20)  (.Q (Ex_D1[20]), .C (CLK_int), .CE (EN_int), .D (
         nx18439z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(19)  (.Q (Ex_D1[19]), .C (CLK_int), .CE (EN_int), .D (
         nx20435z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(18)  (.Q (Ex_D1[18]), .C (CLK_int), .CE (EN_int), .D (
         nx21432z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(17)  (.Q (Ex_D1[17]), .C (CLK_int), .CE (EN_int), .D (
         nx22429z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(16)  (.Q (Ex_D1[16]), .C (CLK_int), .CE (EN_int), .D (
         nx23426z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(15)  (.Q (Ex_D1[15]), .C (CLK_int), .CE (EN_int), .D (
         nx24423z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(14)  (.Q (Ex_D1[14]), .C (CLK_int), .CE (EN_int), .D (
         nx25420z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(13)  (.Q (Ex_D1[13]), .C (CLK_int), .CE (EN_int), .D (
         nx26417z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(12)  (.Q (Ex_D1[12]), .C (CLK_int), .CE (EN_int), .D (
         nx27414z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(11)  (.Q (Ex_D1[11]), .C (CLK_int), .CE (EN_int), .D (
         nx28411z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(10)  (.Q (Ex_D1[10]), .C (CLK_int), .CE (EN_int), .D (
         nx29408z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(9)  (.Q (Ex_D1[9]), .C (CLK_int), .CE (EN_int), .D (
         nx59700z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(8)  (.Q (Ex_D1[8]), .C (CLK_int), .CE (EN_int), .D (
         nx60697z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(7)  (.Q (Ex_D1[7]), .C (CLK_int), .CE (EN_int), .D (
         nx61694z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(6)  (.Q (Ex_D1[6]), .C (CLK_int), .CE (EN_int), .D (
         nx62691z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(5)  (.Q (Ex_D1[5]), .C (CLK_int), .CE (EN_int), .D (
         nx63688z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(4)  (.Q (Ex_D1[4]), .C (CLK_int), .CE (EN_int), .D (
         nx64685z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(3)  (.Q (Ex_D1[3]), .C (CLK_int), .CE (EN_int), .D (nx146z1)
         , .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(2)  (.Q (Ex_D1[2]), .C (CLK_int), .CE (EN_int), .D (nx1143z1
         ), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(1)  (.Q (Ex_D1[1]), .C (CLK_int), .CE (EN_int), .D (nx2140z1
         ), .R (nx59962z2)) ;
    FDRE \reg_Ex_D1(0)  (.Q (Ex_D1[0]), .C (CLK_int), .CE (EN_int), .D (nx3137z1
         ), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(31)  (.Q (Ex_D2[31]), .C (CLK_int), .CE (EN_int), .D (
         nx53928z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(30)  (.Q (Ex_D2[30]), .C (CLK_int), .CE (EN_int), .D (
         nx52931z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(29)  (.Q (Ex_D2[29]), .C (CLK_int), .CE (EN_int), .D (
         nx50935z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(28)  (.Q (Ex_D2[28]), .C (CLK_int), .CE (EN_int), .D (
         nx49938z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(27)  (.Q (Ex_D2[27]), .C (CLK_int), .CE (EN_int), .D (
         nx48941z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(26)  (.Q (Ex_D2[26]), .C (CLK_int), .CE (EN_int), .D (
         nx47944z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(25)  (.Q (Ex_D2[25]), .C (CLK_int), .CE (EN_int), .D (
         nx46947z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(24)  (.Q (Ex_D2[24]), .C (CLK_int), .CE (EN_int), .D (
         nx45950z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(23)  (.Q (Ex_D2[23]), .C (CLK_int), .CE (EN_int), .D (
         nx44953z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(22)  (.Q (Ex_D2[22]), .C (CLK_int), .CE (EN_int), .D (
         nx43956z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(21)  (.Q (Ex_D2[21]), .C (CLK_int), .CE (EN_int), .D (
         nx42959z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(20)  (.Q (Ex_D2[20]), .C (CLK_int), .CE (EN_int), .D (
         nx41962z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(19)  (.Q (Ex_D2[19]), .C (CLK_int), .CE (EN_int), .D (
         nx39966z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(18)  (.Q (Ex_D2[18]), .C (CLK_int), .CE (EN_int), .D (
         nx38969z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(17)  (.Q (Ex_D2[17]), .C (CLK_int), .CE (EN_int), .D (
         nx37972z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(16)  (.Q (Ex_D2[16]), .C (CLK_int), .CE (EN_int), .D (
         nx36975z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(15)  (.Q (Ex_D2[15]), .C (CLK_int), .CE (EN_int), .D (
         nx35978z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(14)  (.Q (Ex_D2[14]), .C (CLK_int), .CE (EN_int), .D (
         nx34981z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(13)  (.Q (Ex_D2[13]), .C (CLK_int), .CE (EN_int), .D (
         nx33984z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(12)  (.Q (Ex_D2[12]), .C (CLK_int), .CE (EN_int), .D (
         nx32987z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(11)  (.Q (Ex_D2[11]), .C (CLK_int), .CE (EN_int), .D (
         nx31990z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(10)  (.Q (Ex_D2[10]), .C (CLK_int), .CE (EN_int), .D (
         nx30993z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(9)  (.Q (Ex_D2[9]), .C (CLK_int), .CE (EN_int), .D (
         nx62953z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(8)  (.Q (Ex_D2[8]), .C (CLK_int), .CE (EN_int), .D (
         nx61956z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(7)  (.Q (Ex_D2[7]), .C (CLK_int), .CE (EN_int), .D (
         nx60959z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(6)  (.Q (Ex_D2[6]), .C (CLK_int), .CE (EN_int), .D (
         nx59962z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(5)  (.Q (Ex_D2[5]), .C (CLK_int), .CE (EN_int), .D (
         nx58965z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(4)  (.Q (Ex_D2[4]), .C (CLK_int), .CE (EN_int), .D (
         nx57968z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(3)  (.Q (Ex_D2[3]), .C (CLK_int), .CE (EN_int), .D (
         nx56971z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(2)  (.Q (Ex_D2[2]), .C (CLK_int), .CE (EN_int), .D (
         nx55974z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(1)  (.Q (Ex_D2[1]), .C (CLK_int), .CE (EN_int), .D (
         nx54977z1), .R (nx59962z2)) ;
    FDRE \reg_Ex_D2(0)  (.Q (Ex_D2[0]), .C (CLK_int), .CE (EN_int), .D (
         nx53980z1), .R (nx59962z2)) ;
    FDRE \reg_Mem_Alu_R(6)  (.Q (Mem_Alu_R[6]), .C (CLK_int), .CE (EN_int), .D (
         nx30553z1), .R (nx58593z1)) ;
    FDRE \reg_Mem_Alu_R(5)  (.Q (Mem_Alu_R[5]), .C (CLK_int), .CE (EN_int), .D (
         nx29556z1), .R (nx58593z1)) ;
    FDRE \reg_Mem_Alu_R(4)  (.Q (Mem_Alu_R[4]), .C (CLK_int), .CE (EN_int), .D (
         nx28559z1), .R (nx58593z1)) ;
    FDRE \reg_Mem_Alu_R(3)  (.Q (Mem_Alu_R[3]), .C (CLK_int), .CE (EN_int), .D (
         nx27562z1), .R (nx58593z1)) ;
    FDRE \reg_Mem_Alu_R(2)  (.Q (Mem_Alu_R[2]), .C (CLK_int), .CE (EN_int), .D (
         nx26565z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(31)  (.Q (Wb_D[31]), .C (CLK_int), .CE (EN_int), .D (nx4630z1
         ), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(30)  (.Q (Wb_D[30]), .C (CLK_int), .CE (EN_int), .D (nx3633z1
         ), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(29)  (.Q (Wb_D[29]), .C (CLK_int), .CE (EN_int), .D (nx1637z1
         ), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(28)  (.Q (Wb_D[28]), .C (CLK_int), .CE (EN_int), .D (nx640z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(27)  (.Q (Wb_D[27]), .C (CLK_int), .CE (EN_int), .D (
         nx65179z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(26)  (.Q (Wb_D[26]), .C (CLK_int), .CE (EN_int), .D (
         nx64182z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(25)  (.Q (Wb_D[25]), .C (CLK_int), .CE (EN_int), .D (
         nx63185z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(24)  (.Q (Wb_D[24]), .C (CLK_int), .CE (EN_int), .D (
         nx62188z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(23)  (.Q (Wb_D[23]), .C (CLK_int), .CE (EN_int), .D (
         nx61191z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(22)  (.Q (Wb_D[22]), .C (CLK_int), .CE (EN_int), .D (
         nx60194z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(21)  (.Q (Wb_D[21]), .C (CLK_int), .CE (EN_int), .D (
         nx59197z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(20)  (.Q (Wb_D[20]), .C (CLK_int), .CE (EN_int), .D (
         nx58200z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(19)  (.Q (Wb_D[19]), .C (CLK_int), .CE (EN_int), .D (
         nx56204z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(18)  (.Q (Wb_D[18]), .C (CLK_int), .CE (EN_int), .D (
         nx55207z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(17)  (.Q (Wb_D[17]), .C (CLK_int), .CE (EN_int), .D (
         nx54210z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(16)  (.Q (Wb_D[16]), .C (CLK_int), .CE (EN_int), .D (
         nx53213z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(15)  (.Q (Wb_D[15]), .C (CLK_int), .CE (EN_int), .D (
         nx52216z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(14)  (.Q (Wb_D[14]), .C (CLK_int), .CE (EN_int), .D (
         nx51219z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(13)  (.Q (Wb_D[13]), .C (CLK_int), .CE (EN_int), .D (
         nx50222z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(12)  (.Q (Wb_D[12]), .C (CLK_int), .CE (EN_int), .D (
         nx49225z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(11)  (.Q (Wb_D[11]), .C (CLK_int), .CE (EN_int), .D (
         nx48228z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(10)  (.Q (Wb_D[10]), .C (CLK_int), .CE (EN_int), .D (
         nx47231z1), .R (nx58593z1)) ;
    FDRE \reg_Wb_D(9)  (.Q (Wb_D[9]), .C (CLK_int), .CE (EN_int), .D (nx7359z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(8)  (.Q (Wb_D[8]), .C (CLK_int), .CE (EN_int), .D (nx6362z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(7)  (.Q (Wb_D[7]), .C (CLK_int), .CE (EN_int), .D (nx5365z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(6)  (.Q (Wb_D[6]), .C (CLK_int), .CE (EN_int), .D (nx4368z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(5)  (.Q (Wb_D[5]), .C (CLK_int), .CE (EN_int), .D (nx3371z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(4)  (.Q (Wb_D[4]), .C (CLK_int), .CE (EN_int), .D (nx2374z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(3)  (.Q (Wb_D[3]), .C (CLK_int), .CE (EN_int), .D (nx1377z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(2)  (.Q (Wb_D[2]), .C (CLK_int), .CE (EN_int), .D (nx380z1), 
         .R (nx58593z1)) ;
    FDRE \reg_Wb_D(1)  (.Q (Wb_D[1]), .C (CLK_int), .CE (EN_int), .D (nx64919z1)
         , .R (nx58593z1)) ;
    FDRE \reg_Wb_D(0)  (.Q (Wb_D[0]), .C (CLK_int), .CE (EN_int), .D (nx63922z1)
         , .R (nx58593z1)) ;
    FDRE \pc_reg_addr(31)  (.Q (Addr_1_0[31]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[31]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(30)  (.Q (Addr_1_0[30]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[30]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(29)  (.Q (Addr_1_0[29]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[29]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(28)  (.Q (Addr_1_0[28]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[28]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(27)  (.Q (Addr_1_0[27]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[27]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(26)  (.Q (Addr_1_0[26]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[26]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(25)  (.Q (Addr_1_0[25]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[25]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(24)  (.Q (Addr_1_0[24]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[24]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(23)  (.Q (Addr_1_0[23]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[23]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(22)  (.Q (Addr_1_0[22]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[22]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(21)  (.Q (Addr_1_0[21]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[21]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(20)  (.Q (Addr_1_0[20]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[20]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(19)  (.Q (Addr_1_0[19]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[19]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(18)  (.Q (Addr_1_0[18]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[18]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(17)  (.Q (Addr_1_0[17]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[17]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(16)  (.Q (Addr_1_0[16]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[16]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(15)  (.Q (Addr_1_0[15]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[15]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(14)  (.Q (Addr_1_0[14]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[14]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(13)  (.Q (Addr_1_0[13]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[13]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(12)  (.Q (Addr_1_0[12]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[12]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(11)  (.Q (Addr_1_0[11]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[11]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(10)  (.Q (Addr_1_0[10]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[10]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(9)  (.Q (Addr_1_0[9]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[9]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(8)  (.Q (Addr_1_0[8]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[8]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(7)  (.Q (Addr_1_0[7]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[7]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(6)  (.Q (Addr_1_0[6]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[6]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(5)  (.Q (Addr_1_0[5]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[5]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(4)  (.Q (Addr_1_0[4]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[4]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(3)  (.Q (Addr_1_0[3]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[3]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(2)  (.Q (Addr_1_0[2]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[2]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(1)  (.Q (Addr_1_0[1]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[1]), .R (pc_not_clr_n)) ;
    FDRE \pc_reg_addr(0)  (.Q (Addr_1_0[0]), .C (CLK_int), .CE (nx42977z1), .D (
         Next_Addr[0]), .R (pc_not_clr_n)) ;
    FDRE \if_id_reg_ID_pc_add4(31)  (.Q (Id_Pc_Add4[31]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(31)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(30)  (.Q (Id_Pc_Add4[30]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(30)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(29)  (.Q (Id_Pc_Add4[29]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(29)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(28)  (.Q (Id_Pc_Add4[28]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(28)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(27)  (.Q (Id_Pc_Add4[27]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(27)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(26)  (.Q (Id_Pc_Add4[26]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(26)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(25)  (.Q (Id_Pc_Add4[25]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(25)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(24)  (.Q (Id_Pc_Add4[24]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(24)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(23)  (.Q (Id_Pc_Add4[23]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(23)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(22)  (.Q (Id_Pc_Add4[22]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(22)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(21)  (.Q (Id_Pc_Add4[21]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(21)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(20)  (.Q (Id_Pc_Add4[20]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(20)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(19)  (.Q (Id_Pc_Add4[19]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(19)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(18)  (.Q (Id_Pc_Add4[18]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(18)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(17)  (.Q (Id_Pc_Add4[17]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(17)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(16)  (.Q (Id_Pc_Add4[16]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(16)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(15)  (.Q (Id_Pc_Add4[15]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(15)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(14)  (.Q (Id_Pc_Add4[14]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(14)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(13)  (.Q (Id_Pc_Add4[13]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(13)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(12)  (.Q (Id_Pc_Add4[12]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(12)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(11)  (.Q (Id_Pc_Add4[11]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(11)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(10)  (.Q (Id_Pc_Add4[10]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(10)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(9)  (.Q (Id_Pc_Add4[9]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(9)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(8)  (.Q (Id_Pc_Add4[8]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(8)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(7)  (.Q (Id_Pc_Add4[7]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(7)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(6)  (.Q (Id_Pc_Add4[6]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(6)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(5)  (.Q (Id_Pc_Add4[5]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(5)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(4)  (.Q (Id_Pc_Add4[4]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(4)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(3)  (.Q (Id_Pc_Add4[3]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(3)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(2)  (.Q (Id_Pc_Add4[2]), .C (CLK_int), .CE (
         nx42977z1), .D (\Pc_Add4(2)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(1)  (.Q (Id_Pc_Add4[1]), .C (CLK_int), .CE (
         nx42977z1), .D (Addr_1_0[1]), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_pc_add4(0)  (.Q (Id_Pc_Add4[0]), .C (CLK_int), .CE (
         nx42977z1), .D (Addr_1_0[0]), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(29)  (.Q (\Id_Inst(29)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(29)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(28)  (.Q (\Id_Inst(28)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(28)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(26)  (.Q (\Id_Inst(26)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(31)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(13)  (.Q (\Id_Extimm(13)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(13)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(12)  (.Q (\Id_Extimm(12)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(12)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(11)  (.Q (\Id_Extimm(11)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(11)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(4)  (.Q (\Id_Extimm(4)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(4)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(3)  (.Q (\Id_Extimm(3)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(3)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(2)  (.Q (\Id_Extimm(2)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(2)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(1)  (.Q (\Id_Extimm(1)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(1)  ), .R (nx28580z1)) ;
    FDRE \if_id_reg_ID_inst(0)  (.Q (\Id_Extimm(0)  ), .C (CLK_int), .CE (
         nx42977z1), .D (\Instruction(0)  ), .R (nx28580z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(31)  (.Q (Wb_Alu_R[31]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[31]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(30)  (.Q (Wb_Alu_R[30]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[30]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(29)  (.Q (Wb_Alu_R[29]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[29]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(28)  (.Q (Wb_Alu_R[28]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[28]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(27)  (.Q (Wb_Alu_R[27]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[27]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(26)  (.Q (Wb_Alu_R[26]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[26]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(25)  (.Q (Wb_Alu_R[25]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[25]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(24)  (.Q (Wb_Alu_R[24]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[24]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(23)  (.Q (Wb_Alu_R[23]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[23]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(22)  (.Q (Wb_Alu_R[22]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[22]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(21)  (.Q (Wb_Alu_R[21]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[21]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(20)  (.Q (Wb_Alu_R[20]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[20]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(19)  (.Q (Wb_Alu_R[19]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[19]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(18)  (.Q (Wb_Alu_R[18]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[18]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(17)  (.Q (Wb_Alu_R[17]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[17]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(16)  (.Q (Wb_Alu_R[16]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[16]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(15)  (.Q (Wb_Alu_R[15]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[15]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(14)  (.Q (Wb_Alu_R[14]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[14]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(13)  (.Q (Wb_Alu_R[13]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[13]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(12)  (.Q (Wb_Alu_R[12]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[12]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(11)  (.Q (Wb_Alu_R[11]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[11]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(10)  (.Q (Wb_Alu_R[10]), .C (CLK_int), .CE (EN_int
         ), .D (Mem_Alu_R[10]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(9)  (.Q (Wb_Alu_R[9]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[9]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(8)  (.Q (Wb_Alu_R[8]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[8]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(7)  (.Q (Wb_Alu_R[7]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[7]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(6)  (.Q (Wb_Alu_R[6]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[6]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(5)  (.Q (Wb_Alu_R[5]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[5]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(4)  (.Q (Wb_Alu_R[4]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[4]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(3)  (.Q (Wb_Alu_R[3]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[3]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(2)  (.Q (Wb_Alu_R[2]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[2]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(1)  (.Q (Wb_Alu_R[1]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[1]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Alu_R(0)  (.Q (Wb_Alu_R[0]), .C (CLK_int), .CE (EN_int)
         , .D (Mem_Alu_R[0]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Rd(2)  (.Q (\Rd_1_0(2)  ), .C (CLK_int), .CE (EN_int), .D (
         Mem_Rd[2]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Rd(1)  (.Q (\Rd_1_0(1)  ), .C (CLK_int), .CE (EN_int), .D (
         Mem_Rd[1]), .R (nx58593z1)) ;
    FDRE \mem_wb_reg_Wb_Rd(0)  (.Q (\Rd_1_0(0)  ), .C (CLK_int), .CE (EN_int), .D (
         Mem_Rd[0]), .R (nx58593z1)) ;
    FDRE mem_wb_reg_Wb_Reg2reg (.Q (Wb_Reg2reg), .C (CLK_int), .CE (EN_int), .D (
         Mem_Reg2reg), .R (nx58593z1)) ;
    FDRE mem_wb_reg_Wb_Wreg (.Q (Wb_Wreg), .C (CLK_int), .CE (EN_int), .D (
         Mem_Wreg), .R (nx58593z1)) ;
    OBUF \Rd_obuf(0)  (.O (Rd[0]), .I (\Rd_1_0(0)  )) ;
    OBUF \Rd_obuf(1)  (.O (Rd[1]), .I (\Rd_1_0(1)  )) ;
    OBUF \Rd_obuf(2)  (.O (Rd[2]), .I (\Rd_1_0(2)  )) ;
    OBUF \Rd_obuf(3)  (.O (Rd[3]), .I (nx57674z45)) ;
    OBUF \Rd_obuf(4)  (.O (Rd[4]), .I (nx57674z45)) ;
    OBUF \Rt_obuf(0)  (.O (Rt[0]), .I (\Rt_1_0(0)  )) ;
    OBUF \Rt_obuf(1)  (.O (Rt[1]), .I (\Rt_1_0(1)  )) ;
    OBUF \Rt_obuf(2)  (.O (Rt[2]), .I (\Rt_1_0(2)  )) ;
    OBUF \Rt_obuf(3)  (.O (Rt[3]), .I (nx57674z45)) ;
    OBUF \Rt_obuf(4)  (.O (Rt[4]), .I (nx57674z45)) ;
    OBUF \Rs_obuf(0)  (.O (Rs[0]), .I (\Rs_1_0(0)  )) ;
    OBUF \Rs_obuf(1)  (.O (Rs[1]), .I (\Rs_1_0(1)  )) ;
    OBUF \Rs_obuf(2)  (.O (Rs[2]), .I (\Rs_1_0(2)  )) ;
    OBUF \Rs_obuf(3)  (.O (Rs[3]), .I (nx57674z45)) ;
    OBUF \Rs_obuf(4)  (.O (Rs[4]), .I (nx57674z45)) ;
    OBUF condition_met_obuf (.O (condition_met), .I (nx4583z1)) ;
    OBUF stall_obuf (.O (stall), .I (nx42977z2)) ;
    OBUF \Write_D_obuf(0)  (.O (Write_D[0]), .I (nx17673z32)) ;
    OBUF \Write_D_obuf(1)  (.O (Write_D[1]), .I (nx17673z31)) ;
    OBUF \Write_D_obuf(2)  (.O (Write_D[2]), .I (nx17673z30)) ;
    OBUF \Write_D_obuf(3)  (.O (Write_D[3]), .I (nx17673z29)) ;
    OBUF \Write_D_obuf(4)  (.O (Write_D[4]), .I (nx17673z28)) ;
    OBUF \Write_D_obuf(5)  (.O (Write_D[5]), .I (nx17673z27)) ;
    OBUF \Write_D_obuf(6)  (.O (Write_D[6]), .I (nx17673z26)) ;
    OBUF \Write_D_obuf(7)  (.O (Write_D[7]), .I (nx17673z25)) ;
    OBUF \Write_D_obuf(8)  (.O (Write_D[8]), .I (nx17673z24)) ;
    OBUF \Write_D_obuf(9)  (.O (Write_D[9]), .I (nx17673z23)) ;
    OBUF \Write_D_obuf(10)  (.O (Write_D[10]), .I (nx17673z22)) ;
    OBUF \Write_D_obuf(11)  (.O (Write_D[11]), .I (nx17673z21)) ;
    OBUF \Write_D_obuf(12)  (.O (Write_D[12]), .I (nx17673z20)) ;
    OBUF \Write_D_obuf(13)  (.O (Write_D[13]), .I (nx17673z19)) ;
    OBUF \Write_D_obuf(14)  (.O (Write_D[14]), .I (nx17673z18)) ;
    OBUF \Write_D_obuf(15)  (.O (Write_D[15]), .I (nx17673z17)) ;
    OBUF \Write_D_obuf(16)  (.O (Write_D[16]), .I (nx17673z16)) ;
    OBUF \Write_D_obuf(17)  (.O (Write_D[17]), .I (nx17673z15)) ;
    OBUF \Write_D_obuf(18)  (.O (Write_D[18]), .I (nx17673z14)) ;
    OBUF \Write_D_obuf(19)  (.O (Write_D[19]), .I (nx17673z13)) ;
    OBUF \Write_D_obuf(20)  (.O (Write_D[20]), .I (nx17673z12)) ;
    OBUF \Write_D_obuf(21)  (.O (Write_D[21]), .I (nx17673z11)) ;
    OBUF \Write_D_obuf(22)  (.O (Write_D[22]), .I (nx17673z10)) ;
    OBUF \Write_D_obuf(23)  (.O (Write_D[23]), .I (nx17673z9)) ;
    OBUF \Write_D_obuf(24)  (.O (Write_D[24]), .I (nx17673z8)) ;
    OBUF \Write_D_obuf(25)  (.O (Write_D[25]), .I (nx17673z7)) ;
    OBUF \Write_D_obuf(26)  (.O (Write_D[26]), .I (nx17673z6)) ;
    OBUF \Write_D_obuf(27)  (.O (Write_D[27]), .I (nx17673z5)) ;
    OBUF \Write_D_obuf(28)  (.O (Write_D[28]), .I (nx17673z4)) ;
    OBUF \Write_D_obuf(29)  (.O (Write_D[29]), .I (nx17673z3)) ;
    OBUF \Write_D_obuf(30)  (.O (Write_D[30]), .I (nx17673z2)) ;
    OBUF \Write_D_obuf(31)  (.O (Write_D[31]), .I (nx17673z1)) ;
    OBUF \Ex_Alu_R_obuf(0)  (.O (Ex_Alu_R[0]), .I (nx54097z51)) ;
    OBUF \Ex_Alu_R_obuf(1)  (.O (Ex_Alu_R[1]), .I (nx54097z52)) ;
    OBUF \Ex_Alu_R_obuf(2)  (.O (Ex_Alu_R[2]), .I (nx26565z1)) ;
    OBUF \Ex_Alu_R_obuf(3)  (.O (Ex_Alu_R[3]), .I (nx27562z1)) ;
    OBUF \Ex_Alu_R_obuf(4)  (.O (Ex_Alu_R[4]), .I (nx28559z1)) ;
    OBUF \Ex_Alu_R_obuf(5)  (.O (Ex_Alu_R[5]), .I (nx29556z1)) ;
    OBUF \Ex_Alu_R_obuf(6)  (.O (Ex_Alu_R[6]), .I (nx30553z1)) ;
    OBUF \Ex_Alu_R_obuf(7)  (.O (Ex_Alu_R[7]), .I (nx54097z53)) ;
    OBUF \Ex_Alu_R_obuf(8)  (.O (Ex_Alu_R[8]), .I (nx54097z54)) ;
    OBUF \Ex_Alu_R_obuf(9)  (.O (Ex_Alu_R[9]), .I (nx54097z55)) ;
    OBUF \Ex_Alu_R_obuf(10)  (.O (Ex_Alu_R[10]), .I (nx54097z56)) ;
    OBUF \Ex_Alu_R_obuf(11)  (.O (Ex_Alu_R[11]), .I (nx54097z57)) ;
    OBUF \Ex_Alu_R_obuf(12)  (.O (Ex_Alu_R[12]), .I (nx54097z58)) ;
    OBUF \Ex_Alu_R_obuf(13)  (.O (Ex_Alu_R[13]), .I (nx54097z59)) ;
    OBUF \Ex_Alu_R_obuf(14)  (.O (Ex_Alu_R[14]), .I (nx54097z60)) ;
    OBUF \Ex_Alu_R_obuf(15)  (.O (Ex_Alu_R[15]), .I (nx54097z61)) ;
    OBUF \Ex_Alu_R_obuf(16)  (.O (Ex_Alu_R[16]), .I (nx54097z62)) ;
    OBUF \Ex_Alu_R_obuf(17)  (.O (Ex_Alu_R[17]), .I (nx54097z63)) ;
    OBUF \Ex_Alu_R_obuf(18)  (.O (Ex_Alu_R[18]), .I (nx54097z64)) ;
    OBUF \Ex_Alu_R_obuf(19)  (.O (Ex_Alu_R[19]), .I (nx54097z65)) ;
    OBUF \Ex_Alu_R_obuf(20)  (.O (Ex_Alu_R[20]), .I (nx54097z66)) ;
    OBUF \Ex_Alu_R_obuf(21)  (.O (Ex_Alu_R[21]), .I (nx54097z67)) ;
    OBUF \Ex_Alu_R_obuf(22)  (.O (Ex_Alu_R[22]), .I (nx54097z68)) ;
    OBUF \Ex_Alu_R_obuf(23)  (.O (Ex_Alu_R[23]), .I (nx54097z69)) ;
    OBUF \Ex_Alu_R_obuf(24)  (.O (Ex_Alu_R[24]), .I (nx54097z70)) ;
    OBUF \Ex_Alu_R_obuf(25)  (.O (Ex_Alu_R[25]), .I (nx54097z71)) ;
    OBUF \Ex_Alu_R_obuf(26)  (.O (Ex_Alu_R[26]), .I (nx54097z72)) ;
    OBUF \Ex_Alu_R_obuf(27)  (.O (Ex_Alu_R[27]), .I (nx54097z73)) ;
    OBUF \Ex_Alu_R_obuf(28)  (.O (Ex_Alu_R[28]), .I (nx54097z74)) ;
    OBUF \Ex_Alu_R_obuf(29)  (.O (Ex_Alu_R[29]), .I (nx54097z75)) ;
    OBUF \Ex_Alu_R_obuf(30)  (.O (Ex_Alu_R[30]), .I (nx54097z76)) ;
    OBUF \Ex_Alu_R_obuf(31)  (.O (Ex_Alu_R[31]), .I (nx54097z77)) ;
    OBUF \Y_obuf(0)  (.O (Y[0]), .I (nx57674z2)) ;
    OBUF \Y_obuf(1)  (.O (Y[1]), .I (nx14570z1)) ;
    OBUF \Y_obuf(2)  (.O (Y[2]), .I (nx13573z1)) ;
    OBUF \Y_obuf(3)  (.O (Y[3]), .I (nx12576z1)) ;
    OBUF \Y_obuf(4)  (.O (Y[4]), .I (nx11579z1)) ;
    OBUF \Y_obuf(5)  (.O (Y[5]), .I (nx10582z1)) ;
    OBUF \Y_obuf(6)  (.O (Y[6]), .I (nx9585z1)) ;
    OBUF \Y_obuf(7)  (.O (Y[7]), .I (nx54097z38)) ;
    OBUF \Y_obuf(8)  (.O (Y[8]), .I (nx54097z37)) ;
    OBUF \Y_obuf(9)  (.O (Y[9]), .I (nx54097z41)) ;
    OBUF \Y_obuf(10)  (.O (Y[10]), .I (nx54097z40)) ;
    OBUF \Y_obuf(11)  (.O (Y[11]), .I (nx34817z1)) ;
    OBUF \Y_obuf(12)  (.O (Y[12]), .I (nx33820z1)) ;
    OBUF \Y_obuf(13)  (.O (Y[13]), .I (nx32823z1)) ;
    OBUF \Y_obuf(14)  (.O (Y[14]), .I (nx54097z44)) ;
    OBUF \Y_obuf(15)  (.O (Y[15]), .I (nx54097z47)) ;
    OBUF \Y_obuf(16)  (.O (Y[16]), .I (nx54097z32)) ;
    OBUF \Y_obuf(17)  (.O (Y[17]), .I (nx54097z39)) ;
    OBUF \Y_obuf(18)  (.O (Y[18]), .I (nx54097z50)) ;
    OBUF \Y_obuf(19)  (.O (Y[19]), .I (nx54097z43)) ;
    OBUF \Y_obuf(20)  (.O (Y[20]), .I (nx54097z46)) ;
    OBUF \Y_obuf(21)  (.O (Y[21]), .I (nx54097z45)) ;
    OBUF \Y_obuf(22)  (.O (Y[22]), .I (nx54097z49)) ;
    OBUF \Y_obuf(23)  (.O (Y[23]), .I (nx21854z1)) ;
    OBUF \Y_obuf(24)  (.O (Y[24]), .I (nx54097z48)) ;
    OBUF \Y_obuf(25)  (.O (Y[25]), .I (nx54097z42)) ;
    OBUF \Y_obuf(26)  (.O (Y[26]), .I (nx54097z36)) ;
    OBUF \Y_obuf(27)  (.O (Y[27]), .I (nx54097z35)) ;
    OBUF \Y_obuf(28)  (.O (Y[28]), .I (nx54097z34)) ;
    OBUF \Y_obuf(29)  (.O (Y[29]), .I (nx54097z33)) ;
    OBUF \Y_obuf(30)  (.O (Y[30]), .I (nx54097z31)) ;
    OBUF \Y_obuf(31)  (.O (Y[31]), .I (nx54097z30)) ;
    OBUF \Alu_D1_obuf(0)  (.O (Alu_D1[0]), .I (nx22138z1)) ;
    OBUF \Alu_D1_obuf(1)  (.O (Alu_D1[1]), .I (nx21141z1)) ;
    OBUF \Alu_D1_obuf(2)  (.O (Alu_D1[2]), .I (nx20144z1)) ;
    OBUF \Alu_D1_obuf(3)  (.O (Alu_D1[3]), .I (nx19147z1)) ;
    OBUF \Alu_D1_obuf(4)  (.O (Alu_D1[4]), .I (nx18150z1)) ;
    OBUF \Alu_D1_obuf(5)  (.O (Alu_D1[5]), .I (nx17153z1)) ;
    OBUF \Alu_D1_obuf(6)  (.O (Alu_D1[6]), .I (nx16156z1)) ;
    OBUF \Alu_D1_obuf(7)  (.O (Alu_D1[7]), .I (nx15159z1)) ;
    OBUF \Alu_D1_obuf(8)  (.O (Alu_D1[8]), .I (nx14162z1)) ;
    OBUF \Alu_D1_obuf(9)  (.O (Alu_D1[9]), .I (nx13165z1)) ;
    OBUF \Alu_D1_obuf(10)  (.O (Alu_D1[10]), .I (nx33501z1)) ;
    OBUF \Alu_D1_obuf(11)  (.O (Alu_D1[11]), .I (nx32504z1)) ;
    OBUF \Alu_D1_obuf(12)  (.O (Alu_D1[12]), .I (nx31507z1)) ;
    OBUF \Alu_D1_obuf(13)  (.O (Alu_D1[13]), .I (nx30510z1)) ;
    OBUF \Alu_D1_obuf(14)  (.O (Alu_D1[14]), .I (nx29513z1)) ;
    OBUF \Alu_D1_obuf(15)  (.O (Alu_D1[15]), .I (nx28516z1)) ;
    OBUF \Alu_D1_obuf(16)  (.O (Alu_D1[16]), .I (nx27519z1)) ;
    OBUF \Alu_D1_obuf(17)  (.O (Alu_D1[17]), .I (nx26522z1)) ;
    OBUF \Alu_D1_obuf(18)  (.O (Alu_D1[18]), .I (nx25525z1)) ;
    OBUF \Alu_D1_obuf(19)  (.O (Alu_D1[19]), .I (nx24528z1)) ;
    OBUF \Alu_D1_obuf(20)  (.O (Alu_D1[20]), .I (nx22532z1)) ;
    OBUF \Alu_D1_obuf(21)  (.O (Alu_D1[21]), .I (nx21535z1)) ;
    OBUF \Alu_D1_obuf(22)  (.O (Alu_D1[22]), .I (nx20538z1)) ;
    OBUF \Alu_D1_obuf(23)  (.O (Alu_D1[23]), .I (nx19541z1)) ;
    OBUF \Alu_D1_obuf(24)  (.O (Alu_D1[24]), .I (nx18544z1)) ;
    OBUF \Alu_D1_obuf(25)  (.O (Alu_D1[25]), .I (nx17547z1)) ;
    OBUF \Alu_D1_obuf(26)  (.O (Alu_D1[26]), .I (nx16550z1)) ;
    OBUF \Alu_D1_obuf(27)  (.O (Alu_D1[27]), .I (nx15553z1)) ;
    OBUF \Alu_D1_obuf(28)  (.O (Alu_D1[28]), .I (nx14556z1)) ;
    OBUF \Alu_D1_obuf(29)  (.O (Alu_D1[29]), .I (nx13559z1)) ;
    OBUF \Alu_D1_obuf(30)  (.O (Alu_D1[30]), .I (nx11563z1)) ;
    OBUF \Alu_D1_obuf(31)  (.O (Alu_D1[31]), .I (nx10566z1)) ;
    OBUF \Addr_obuf(0)  (.O (Addr[0]), .I (Addr_1_0[0])) ;
    OBUF \Addr_obuf(1)  (.O (Addr[1]), .I (Addr_1_0[1])) ;
    OBUF \Addr_obuf(2)  (.O (Addr[2]), .I (Addr_1_0[2])) ;
    OBUF \Addr_obuf(3)  (.O (Addr[3]), .I (Addr_1_0[3])) ;
    OBUF \Addr_obuf(4)  (.O (Addr[4]), .I (Addr_1_0[4])) ;
    OBUF \Addr_obuf(5)  (.O (Addr[5]), .I (Addr_1_0[5])) ;
    OBUF \Addr_obuf(6)  (.O (Addr[6]), .I (Addr_1_0[6])) ;
    OBUF \Addr_obuf(7)  (.O (Addr[7]), .I (Addr_1_0[7])) ;
    OBUF \Addr_obuf(8)  (.O (Addr[8]), .I (Addr_1_0[8])) ;
    OBUF \Addr_obuf(9)  (.O (Addr[9]), .I (Addr_1_0[9])) ;
    OBUF \Addr_obuf(10)  (.O (Addr[10]), .I (Addr_1_0[10])) ;
    OBUF \Addr_obuf(11)  (.O (Addr[11]), .I (Addr_1_0[11])) ;
    OBUF \Addr_obuf(12)  (.O (Addr[12]), .I (Addr_1_0[12])) ;
    OBUF \Addr_obuf(13)  (.O (Addr[13]), .I (Addr_1_0[13])) ;
    OBUF \Addr_obuf(14)  (.O (Addr[14]), .I (Addr_1_0[14])) ;
    OBUF \Addr_obuf(15)  (.O (Addr[15]), .I (Addr_1_0[15])) ;
    OBUF \Addr_obuf(16)  (.O (Addr[16]), .I (Addr_1_0[16])) ;
    OBUF \Addr_obuf(17)  (.O (Addr[17]), .I (Addr_1_0[17])) ;
    OBUF \Addr_obuf(18)  (.O (Addr[18]), .I (Addr_1_0[18])) ;
    OBUF \Addr_obuf(19)  (.O (Addr[19]), .I (Addr_1_0[19])) ;
    OBUF \Addr_obuf(20)  (.O (Addr[20]), .I (Addr_1_0[20])) ;
    OBUF \Addr_obuf(21)  (.O (Addr[21]), .I (Addr_1_0[21])) ;
    OBUF \Addr_obuf(22)  (.O (Addr[22]), .I (Addr_1_0[22])) ;
    OBUF \Addr_obuf(23)  (.O (Addr[23]), .I (Addr_1_0[23])) ;
    OBUF \Addr_obuf(24)  (.O (Addr[24]), .I (Addr_1_0[24])) ;
    OBUF \Addr_obuf(25)  (.O (Addr[25]), .I (Addr_1_0[25])) ;
    OBUF \Addr_obuf(26)  (.O (Addr[26]), .I (Addr_1_0[26])) ;
    OBUF \Addr_obuf(27)  (.O (Addr[27]), .I (Addr_1_0[27])) ;
    OBUF \Addr_obuf(28)  (.O (Addr[28]), .I (Addr_1_0[28])) ;
    OBUF \Addr_obuf(29)  (.O (Addr[29]), .I (Addr_1_0[29])) ;
    OBUF \Addr_obuf(30)  (.O (Addr[30]), .I (Addr_1_0[30])) ;
    OBUF \Addr_obuf(31)  (.O (Addr[31]), .I (Addr_1_0[31])) ;
    IBUF CLR_N_ibuf (.O (CLR_N_int), .I (CLR_N)) ;
    IBUF EN_ibuf (.O (EN_int), .I (EN)) ;
    VCC ps_vcc (.P (nx15902z32)) ;
    GND ps_gnd (.G (nx57674z45)) ;
    (* HLUTNM = "LUT62_7_16" *)
    LUT3 ix17673z1547 (.O (nx17673z32), .I0 (Wb_D[0]), .I1 (Wb_Alu_R[0]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1547.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_16" *)
    LUT3 ix17673z1546 (.O (nx17673z31), .I0 (Wb_D[1]), .I1 (Wb_Alu_R[1]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1546.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_15" *)
    LUT3 ix17673z1545 (.O (nx17673z30), .I0 (Wb_D[2]), .I1 (Wb_Alu_R[2]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1545.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_15" *)
    LUT3 ix17673z1544 (.O (nx17673z29), .I0 (Wb_D[3]), .I1 (Wb_Alu_R[3]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1544.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_14" *)
    LUT3 ix17673z1543 (.O (nx17673z28), .I0 (Wb_D[4]), .I1 (Wb_Alu_R[4]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1543.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_14" *)
    LUT3 ix17673z1542 (.O (nx17673z27), .I0 (Wb_D[5]), .I1 (Wb_Alu_R[5]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1542.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_13" *)
    LUT3 ix17673z1541 (.O (nx17673z26), .I0 (Wb_D[6]), .I1 (Wb_Alu_R[6]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1541.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_13" *)
    LUT3 ix17673z1540 (.O (nx17673z25), .I0 (Wb_D[7]), .I1 (Wb_Alu_R[7]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1540.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_12" *)
    LUT3 ix17673z1539 (.O (nx17673z24), .I0 (Wb_D[8]), .I1 (Wb_Alu_R[8]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1539.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_12" *)
    LUT3 ix17673z1538 (.O (nx17673z23), .I0 (Wb_D[9]), .I1 (Wb_Alu_R[9]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1538.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_11" *)
    LUT3 ix17673z1537 (.O (nx17673z22), .I0 (Wb_D[10]), .I1 (Wb_Alu_R[10]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1537.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_11" *)
    LUT3 ix17673z1536 (.O (nx17673z21), .I0 (Wb_D[11]), .I1 (Wb_Alu_R[11]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1536.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_10" *)
    LUT3 ix17673z1535 (.O (nx17673z20), .I0 (Wb_D[12]), .I1 (Wb_Alu_R[12]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1535.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_10" *)
    LUT3 ix17673z1534 (.O (nx17673z19), .I0 (Wb_D[13]), .I1 (Wb_Alu_R[13]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1534.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_9" *)
    LUT3 ix17673z1533 (.O (nx17673z18), .I0 (Wb_D[14]), .I1 (Wb_Alu_R[14]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1533.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_9" *)
    LUT3 ix17673z1532 (.O (nx17673z17), .I0 (Wb_D[15]), .I1 (Wb_Alu_R[15]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1532.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_8" *)
    LUT3 ix17673z1531 (.O (nx17673z16), .I0 (Wb_D[16]), .I1 (Wb_Alu_R[16]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1531.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_8" *)
    LUT3 ix17673z1530 (.O (nx17673z15), .I0 (Wb_D[17]), .I1 (Wb_Alu_R[17]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1530.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_7" *)
    LUT3 ix17673z1529 (.O (nx17673z14), .I0 (Wb_D[18]), .I1 (Wb_Alu_R[18]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1529.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_7" *)
    LUT3 ix17673z1528 (.O (nx17673z13), .I0 (Wb_D[19]), .I1 (Wb_Alu_R[19]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1528.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_6" *)
    LUT3 ix17673z1527 (.O (nx17673z12), .I0 (Wb_D[20]), .I1 (Wb_Alu_R[20]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1527.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_6" *)
    LUT3 ix17673z1526 (.O (nx17673z11), .I0 (Wb_D[21]), .I1 (Wb_Alu_R[21]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1526.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_5" *)
    LUT3 ix17673z1525 (.O (nx17673z10), .I0 (Wb_D[22]), .I1 (Wb_Alu_R[22]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1525.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_5" *)
    LUT3 ix17673z1524 (.O (nx17673z9), .I0 (Wb_D[23]), .I1 (Wb_Alu_R[23]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1524.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_4" *)
    LUT3 ix17673z1523 (.O (nx17673z8), .I0 (Wb_D[24]), .I1 (Wb_Alu_R[24]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1523.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_4" *)
    LUT3 ix17673z1522 (.O (nx17673z7), .I0 (Wb_D[25]), .I1 (Wb_Alu_R[25]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1522.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_3" *)
    LUT3 ix17673z1521 (.O (nx17673z6), .I0 (Wb_D[26]), .I1 (Wb_Alu_R[26]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1521.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_3" *)
    LUT3 ix17673z1520 (.O (nx17673z5), .I0 (Wb_D[27]), .I1 (Wb_Alu_R[27]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1520.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_2" *)
    LUT3 ix17673z1519 (.O (nx17673z4), .I0 (Wb_D[28]), .I1 (Wb_Alu_R[28]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1519.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_2" *)
    LUT3 ix17673z1518 (.O (nx17673z3), .I0 (Wb_D[29]), .I1 (Wb_Alu_R[29]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1518.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_1" *)
    LUT3 ix17673z1517 (.O (nx17673z2), .I0 (Wb_D[30]), .I1 (Wb_Alu_R[30]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1517.INIT = 8'hCA;
    (* HLUTNM = "LUT62_7_1" *)
    LUT3 ix17673z1516 (.O (nx17673z1), .I0 (Wb_D[31]), .I1 (Wb_Alu_R[31]), .I2 (
         Wb_Reg2reg)) ;
         defparam ix17673z1516.INIT = 8'hCA;
    LUT6 ix759z1827 (.O (nx759z65), .I0 (\Rt_1_0(2)  ), .I1 (\Rt_1_0(1)  ), .I2 (
         \Rt_1_0(0)  ), .I3 (\Rd_1_0(2)  ), .I4 (\Rd_1_0(1)  ), .I5 (\Rd_1_0(0)  
         )) ;
         defparam ix759z1827.INIT = 64'h8040201008040200;
    LUT6 ix759z1826 (.O (nx759z32), .I0 (\Rs_1_0(2)  ), .I1 (\Rs_1_0(1)  ), .I2 (
         \Rs_1_0(0)  ), .I3 (\Rd_1_0(2)  ), .I4 (\Rd_1_0(1)  ), .I5 (\Rd_1_0(0)  
         )) ;
         defparam ix759z1826.INIT = 64'h8040201008040200;
    LUT2 ix42977z1318 (.O (nx42977z1), .I0 (nx42977z2), .I1 (EN_int)) ;
         defparam ix42977z1318.INIT = 4'h4;
    LUT2 ix17673z1354 (.O (nx17673z33), .I0 (Wb_Wreg), .I1 (CLR_N_int)) ;
         defparam ix17673z1354.INIT = 4'h8;
    MUX4X32_0 mux4x_32 (.px2900 (nx15902z1), .p_nbus_Next_Addr ({Next_Addr[0],
              Next_Addr[1],Next_Addr[2],Next_Addr[3],Next_Addr[4],Next_Addr[5],
              Next_Addr[6],Next_Addr[7],Next_Addr[8],Next_Addr[9],Next_Addr[10],
              Next_Addr[11],Next_Addr[12],Next_Addr[13],Next_Addr[14],
              Next_Addr[15],Next_Addr[16],Next_Addr[17],Next_Addr[18],
              Next_Addr[19],Next_Addr[20],Next_Addr[21],Next_Addr[22],
              Next_Addr[23],Next_Addr[24],Next_Addr[25],Next_Addr[26],
              Next_Addr[27],Next_Addr[28],Next_Addr[29],Next_Addr[30],
              Next_Addr[31]}), .px2902 (nx15902z2), .px2904 (nx15902z3), .px2906 (
              nx15902z4), .px2908 (nx15902z5), .px2910 (nx15902z6), .px2912 (
              nx15902z7), .px2914 (nx15902z8), .px2916 (nx15902z9), .px2918 (
              nx15902z10), .px2920 (nx15902z11), .px2922 (nx15902z12), .px2924 (
              nx15902z13), .px2926 (nx15902z14), .px2928 (nx15902z15), .px2930 (
              nx15902z16), .px2932 (nx15902z17), .px2934 (nx15902z18), .px2936 (
              nx15902z19), .px2938 (nx15902z20), .px2940 (nx15902z21), .px2942 (
              nx15902z22), .px2944 (nx15902z23), .px2946 (nx15902z24), .px2948 (
              nx15902z25), .px2950 (nx15902z26), .px2952 (nx15902z27), .px2954 (
              nx15902z28), .px2956 (nx15902z29), .px2958 (nx15902z30), .px2960 (
              nx15902z31), .px2855 (nx15902z32), .px2962 (nx15902z33)) ;
    INST_MEM_0 instuction_mem (.p_nbus_Addr_1_0 ({Addr_1_0[9],Addr_1_0[29],
               Addr_1_0[30],Addr_1_0[31],Addr_1_0[25],Addr_1_0[26],Addr_1_0[27],
               Addr_1_0[28],Addr_1_0[17],Addr_1_0[21],Addr_1_0[22],Addr_1_0[24],
               Addr_1_0[18],Addr_1_0[19],Addr_1_0[20],Addr_1_0[23],Addr_1_0[0],
               Addr_1_0[1],Addr_1_0[7],Addr_1_0[8],Addr_1_0[10],Addr_1_0[11],
               Addr_1_0[12],Addr_1_0[16],Addr_1_0[13],Addr_1_0[14],Addr_1_0[15],
               Addr_1_0[2],Addr_1_0[3],Addr_1_0[4],Addr_1_0[5],Addr_1_0[6]}), .\p_Instruction(0)   (
               \Instruction(0)  ), .\p_Instruction(1)   (\Instruction(1)  ), .\p_Instruction(2)   (
               \Instruction(2)  ), .\p_Instruction(3)   (\Instruction(3)  ), .\p_Instruction(4)   (
               \Instruction(4)  ), .\p_Instruction(13)   (\Instruction(13)  ), .\p_Instruction(31)   (
               \Instruction(31)  ), .\p_Instruction(11)   (\Instruction(11)  ), 
               .\p_Instruction(12)   (\Instruction(12)  ), .\p_Instruction(16)   (
               \Instruction(16)  ), .\p_Instruction(17)   (\Instruction(17)  ), 
               .\p_Instruction(18)   (\Instruction(18)  ), .\p_Instruction(21)   (
               \Instruction(21)  ), .\p_Instruction(22)   (\Instruction(22)  ), 
               .\p_Instruction(23)   (\Instruction(23)  ), .\p_Instruction(28)   (
               \Instruction(28)  ), .\p_Instruction(29)   (\Instruction(29)  )
               ) ;
    REG_FILE_unfolded0_0 reg_file (.\p_Rs_1_0(0)   (\Rs_1_0(0)  ), .\p_Rs_1_0(1)   (
                         \Rs_1_0(1)  ), .\p_Rs_1_0(2)   (\Rs_1_0(2)  ), .\p_Rt_1_0(0)   (
                         \Rt_1_0(0)  ), .\p_Rt_1_0(1)   (\Rt_1_0(1)  ), .\p_Rt_1_0(2)   (
                         \Rt_1_0(2)  ), .p_CLR_N_int (CLR_N_int), .\p_Rd_1_0(0)   (
                         \Rd_1_0(0)  ), .\p_Rd_1_0(1)   (\Rd_1_0(1)  ), .\p_Rd_1_0(2)   (
                         \Rd_1_0(2)  ), .p_rtlcs104 (nx759z1), .px3105 (nx6473z1
                         ), .p_rtlcs103 (nx759z2), .px3104 (nx7470z1), .p_rtlcs102 (
                         nx759z3), .px3103 (nx9466z1), .p_rtlcs101 (nx759z4), .px3102 (
                         nx10463z1), .p_rtlcs100 (nx759z5), .px3101 (nx11460z1)
                         , .p_rtlcs99 (nx759z6), .px3100 (nx12457z1), .p_rtlcs98 (
                         nx759z7), .px3099 (nx13454z1), .p_rtlcs97 (nx759z8), .px3098 (
                         nx14451z1), .p_rtlcs96 (nx759z9), .px3097 (nx15448z1), 
                         .p_rtlcs95 (nx759z10), .px3096 (nx16445z1), .p_rtlcs94 (
                         nx759z11), .px3095 (nx17442z1), .p_rtlcs93 (nx759z12), 
                         .px3094 (nx18439z1), .p_rtlcs92 (nx759z13), .px3093 (
                         nx20435z1), .p_rtlcs91 (nx759z14), .px3092 (nx21432z1)
                         , .p_rtlcs90 (nx759z15), .px3091 (nx22429z1), .p_rtlcs89 (
                         nx759z16), .px3090 (nx23426z1), .p_rtlcs88 (nx759z17), 
                         .px3089 (nx24423z1), .p_rtlcs87 (nx759z18), .px3088 (
                         nx25420z1), .p_rtlcs86 (nx759z19), .px3087 (nx26417z1)
                         , .p_rtlcs85 (nx759z20), .px3086 (nx27414z1), .p_rtlcs84 (
                         nx759z21), .px3085 (nx28411z1), .p_rtlcs83 (nx759z22), 
                         .px3084 (nx29408z1), .p_rtlcs82 (nx759z23), .px3083 (
                         nx59700z1), .p_rtlcs81 (nx759z24), .px3082 (nx60697z1)
                         , .p_rtlcs80 (nx759z25), .px3081 (nx61694z1), .p_rtlcs79 (
                         nx759z26), .px3080 (nx62691z1), .p_rtlcs78 (nx759z27), 
                         .px3079 (nx63688z1), .p_rtlcs77 (nx759z28), .px3078 (
                         nx64685z1), .p_rtlcs76 (nx759z29), .px3077 (nx146z1), .p_rtlcs75 (
                         nx759z30), .px3076 (nx1143z1), .p_rtlcs74 (nx759z31), .px3075 (
                         nx2140z1), .px3448 (nx759z32), .p_rtlcs73 (nx759z33), .px3074 (
                         nx3137z1), .p_rtlcs141 (nx759z34), .p_nbus_Wb_Alu_R ({
                         Wb_Alu_R[31],Wb_Alu_R[30],Wb_Alu_R[29],Wb_Alu_R[28],
                         Wb_Alu_R[27],Wb_Alu_R[26],Wb_Alu_R[25],Wb_Alu_R[24],
                         Wb_Alu_R[23],Wb_Alu_R[22],Wb_Alu_R[21],Wb_Alu_R[20],
                         Wb_Alu_R[19],Wb_Alu_R[18],Wb_Alu_R[17],Wb_Alu_R[16],
                         Wb_Alu_R[15],Wb_Alu_R[14],Wb_Alu_R[13],Wb_Alu_R[12],
                         Wb_Alu_R[11],Wb_Alu_R[10],Wb_Alu_R[9],Wb_Alu_R[8],
                         Wb_Alu_R[7],Wb_Alu_R[6],Wb_Alu_R[5],Wb_Alu_R[4],
                         Wb_Alu_R[3],Wb_Alu_R[2],Wb_Alu_R[1],Wb_Alu_R[0]}), .p_nbus_Wb_D (
                         {Wb_D[31],Wb_D[30],Wb_D[29],Wb_D[28],Wb_D[27],Wb_D[26],
                         Wb_D[25],Wb_D[24],Wb_D[23],Wb_D[22],Wb_D[21],Wb_D[20],
                         Wb_D[19],Wb_D[18],Wb_D[17],Wb_D[16],Wb_D[15],Wb_D[14],
                         Wb_D[13],Wb_D[12],Wb_D[11],Wb_D[10],Wb_D[9],Wb_D[8],
                         Wb_D[7],Wb_D[6],Wb_D[5],Wb_D[4],Wb_D[3],Wb_D[2],Wb_D[1]
                         ,Wb_D[0]}), .px3073 (nx53928z1), .p_rtlcs140 (nx759z35)
                         , .px3072 (nx52931z1), .p_rtlcs139 (nx759z36), .px3071 (
                         nx50935z1), .p_rtlcs138 (nx759z37), .px3070 (nx49938z1)
                         , .p_rtlcs137 (nx759z38), .px3069 (nx48941z1), .p_rtlcs136 (
                         nx759z39), .px3068 (nx47944z1), .p_rtlcs135 (nx759z40)
                         , .px3067 (nx46947z1), .p_rtlcs134 (nx759z41), .px3066 (
                         nx45950z1), .p_rtlcs133 (nx759z42), .px3065 (nx44953z1)
                         , .p_rtlcs132 (nx759z43), .px3064 (nx43956z1), .p_rtlcs131 (
                         nx759z44), .px3063 (nx42959z1), .p_rtlcs130 (nx759z45)
                         , .px3062 (nx41962z1), .p_rtlcs129 (nx759z46), .px3061 (
                         nx39966z1), .p_rtlcs128 (nx759z47), .px3060 (nx38969z1)
                         , .p_rtlcs127 (nx759z48), .px3059 (nx37972z1), .p_rtlcs126 (
                         nx759z49), .px3058 (nx36975z1), .p_rtlcs125 (nx759z50)
                         , .px3057 (nx35978z1), .p_rtlcs124 (nx759z51), .px3056 (
                         nx34981z1), .p_rtlcs123 (nx759z52), .px3055 (nx33984z1)
                         , .p_rtlcs122 (nx759z53), .px3054 (nx32987z1), .p_rtlcs121 (
                         nx759z54), .px3053 (nx31990z1), .p_rtlcs120 (nx759z55)
                         , .px3052 (nx30993z1), .p_rtlcs119 (nx759z56), .px3051 (
                         nx62953z1), .p_rtlcs118 (nx759z57), .px3050 (nx61956z1)
                         , .p_rtlcs117 (nx759z58), .px3049 (nx60959z1), .p_rtlcs116 (
                         nx759z59), .px3048 (nx59962z1), .p_rtlcs115 (nx759z60)
                         , .px3047 (nx58965z1), .p_rtlcs114 (nx759z61), .px3046 (
                         nx57968z1), .p_rtlcs113 (nx759z62), .px3045 (nx56971z1)
                         , .p_rtlcs112 (nx759z63), .px3044 (nx55974z1), .p_rtlcs111 (
                         nx759z64), .px3043 (nx54977z1), .px3443 (nx759z65), .p_rtlcs110 (
                         nx759z66), .p_Wb_Reg2reg (Wb_Reg2reg), .px3042 (
                         nx53980z1), .p_pc_not_clr_n (pc_not_clr_n), .p_Wb_Wreg (
                         Wb_Wreg), .p_CLK_int (CLK_int)) ;
    ID_EX_unfolded0_0 id_ex (.\p_Rs_1_0(0)   (\Rs_1_0(0)  ), .\p_Rs_1_0(1)   (
                      \Rs_1_0(1)  ), .\p_Rs_1_0(2)   (\Rs_1_0(2)  ), .px3449 (
                      nx28580z1), .p_CLR_N_int (CLR_N_int), .px3450 (nx4583z1), 
                      .px3452 (nx42977z2), .px3419 (nx57674z32), .px3370 (
                      nx23941z1), .px3371 (nx23941z2), .px3369 (nx57674z2), .px3366 (
                      nx57674z31), .px3350 (nx57674z35), .px3346 (nx57674z36), .px3422 (
                      nx23941z3), .px3423 (nx57674z33), .px3426 (nx23941z4), .px3427 (
                      nx57674z34), .px3430 (nx23941z5), .px3431 (nx23941z6), .px3206 (
                      nx57674z37), .px3367 (nx23941z7), .p_nbus_Ex_D2 ({Ex_D2[1]
                      ,Ex_D2[2],Ex_D2[3],Ex_D2[4],Ex_D2[11],Ex_D2[12]}), .px3003 (
                      nx14570z1), .px3420 (nx23941z8), .px3002 (nx13573z1), .px3424 (
                      nx23941z9), .px3001 (nx12576z1), .px3428 (nx23941z10), .px3000 (
                      nx11579z1), .p_nbus_Mem_Alu_R ({Mem_Alu_R[5],Mem_Alu_R[13]
                      }), .px3432 (nx23941z11), .px2999 (nx10582z1), .px3439 (
                      nx23941z12), .px3462 (nx23941z13), .px2998 (nx9585z1), .px3351 (
                      nx23941z14), .px2997 (nx34817z1), .px3347 (nx23941z15), .px2996 (
                      nx33820z1), .px3343 (nx23941z16), .px2995 (nx32823z1), .\p_Pc_Add4(31)   (
                      \Pc_Add4(31)  ), .px2962 (nx15902z33), .\p_Pc_Add4(30)   (
                      \Pc_Add4(30)  ), .px2960 (nx15902z31), .\p_Pc_Add4(29)   (
                      \Pc_Add4(29)  ), .px2958 (nx15902z30), .\p_Pc_Add4(28)   (
                      \Pc_Add4(28)  ), .px2956 (nx15902z29), .\p_Pc_Add4(27)   (
                      \Pc_Add4(27)  ), .px2954 (nx15902z28), .\p_Pc_Add4(26)   (
                      \Pc_Add4(26)  ), .px2952 (nx15902z27), .\p_Pc_Add4(25)   (
                      \Pc_Add4(25)  ), .px2950 (nx15902z26), .\p_Pc_Add4(24)   (
                      \Pc_Add4(24)  ), .px2948 (nx15902z25), .\p_Pc_Add4(23)   (
                      \Pc_Add4(23)  ), .px2946 (nx15902z24), .\p_Pc_Add4(22)   (
                      \Pc_Add4(22)  ), .px2944 (nx15902z23), .\p_Pc_Add4(21)   (
                      \Pc_Add4(21)  ), .px2942 (nx15902z22), .\p_Pc_Add4(20)   (
                      \Pc_Add4(20)  ), .px2940 (nx15902z21), .\p_Pc_Add4(19)   (
                      \Pc_Add4(19)  ), .px2938 (nx15902z20), .\p_Pc_Add4(18)   (
                      \Pc_Add4(18)  ), .px2936 (nx15902z19), .\p_Pc_Add4(17)   (
                      \Pc_Add4(17)  ), .px2934 (nx15902z18), .\p_Pc_Add4(16)   (
                      \Pc_Add4(16)  ), .px2932 (nx15902z17), .\p_Pc_Add4(15)   (
                      \Pc_Add4(15)  ), .px2930 (nx15902z16), .\p_Pc_Add4(14)   (
                      \Pc_Add4(14)  ), .px2928 (nx15902z15), .\p_Pc_Add4(13)   (
                      \Pc_Add4(13)  ), .px2926 (nx15902z14), .\p_Pc_Add4(12)   (
                      \Pc_Add4(12)  ), .px2924 (nx15902z13), .\p_Pc_Add4(11)   (
                      \Pc_Add4(11)  ), .px2922 (nx15902z12), .\p_Pc_Add4(10)   (
                      \Pc_Add4(10)  ), .px2920 (nx15902z11), .\p_Pc_Add4(9)   (
                      \Pc_Add4(9)  ), .px2918 (nx15902z10), .\p_Pc_Add4(8)   (
                      \Pc_Add4(8)  ), .px2916 (nx15902z9), .\p_Pc_Add4(7)   (
                      \Pc_Add4(7)  ), .px2914 (nx15902z8), .\p_Pc_Add4(6)   (
                      \Pc_Add4(6)  ), .px2912 (nx15902z7), .\p_Pc_Add4(5)   (
                      \Pc_Add4(5)  ), .px2910 (nx15902z6), .\p_Pc_Add4(4)   (
                      \Pc_Add4(4)  ), .px2908 (nx15902z5), .\p_Pc_Add4(3)   (
                      \Pc_Add4(3)  ), .px2906 (nx15902z4), .\p_Pc_Add4(2)   (
                      \Pc_Add4(2)  ), .px2904 (nx15902z3), .p_nbus_Addr_1_0 ({
                      Addr_1_0[1],Addr_1_0[0]}), .px2902 (nx15902z2), .p_Ex_Z (
                      Ex_Z), .px2900 (nx15902z1), .\p_Rt_1_0(2)   (\Rt_1_0(2)  )
                      , .\p_Rt_1_0(1)   (\Rt_1_0(1)  ), .\p_Rt_1_0(0)   (
                      \Rt_1_0(0)  ), .\p_Id_Extimm(0)   (\Id_Extimm(0)  ), .\p_Ex_Extimm(0)   (
                      \Ex_Extimm(0)  ), .\p_Id_Extimm(1)   (\Id_Extimm(1)  ), .\p_Id_Extimm(2)   (
                      \Id_Extimm(2)  ), .\p_Id_Extimm(3)   (\Id_Extimm(3)  ), .\p_Id_Extimm(4)   (
                      \Id_Extimm(4)  ), .\p_Id_Extimm(13)   (\Id_Extimm(13)  ), 
                      .\p_Ex_Extimm(13)   (\Ex_Extimm(13)  ), .\p_Id_Inst(26)   (
                      \Id_Inst(26)  ), .\p_Ex_Op(0)   (\Ex_Op(0)  ), .\p_Id_Extimm(11)   (
                      \Id_Extimm(11)  ), .\p_Id_Extimm(12)   (\Id_Extimm(12)  )
                      , .\p_Id_Inst(28)   (\Id_Inst(28)  ), .\p_Id_Inst(29)   (
                      \Id_Inst(29)  ), .p_nbus_Ex_Rd ({Ex_Rd[0],Ex_Rd[1],
                      Ex_Rd[2]}), .p_nbus_Ex_Aluc ({Ex_Aluc[0],Ex_Aluc[1],
                      Ex_Aluc[2]}), .px3253 (nx23941z17), .p_nbus_Ex_Fwd_A ({
                      Ex_Fwd_A[0],Ex_Fwd_A[1]}), .px3255 (nx54097z29), .px3256 (
                      nx23941z18), .p_nbus_Ex_Fwd_B ({Ex_Fwd_B[0],Ex_Fwd_B[1]})
                      , .px3258 (nx54097z28), .p_Ex_Wreg (Ex_Wreg), .p_Ex_Reg2reg (
                      Ex_Reg2reg), .p_Ex_Wmem (Ex_Wmem), .p_Ex_Aluqb (Ex_Aluqb)
                      , .p_nbus_Id_Pc_Add4 ({Id_Pc_Add4[0],Id_Pc_Add4[1],
                      Id_Pc_Add4[31],Id_Pc_Add4[30],Id_Pc_Add4[29],
                      Id_Pc_Add4[28],Id_Pc_Add4[27],Id_Pc_Add4[26],
                      Id_Pc_Add4[25],Id_Pc_Add4[24],Id_Pc_Add4[23],
                      Id_Pc_Add4[22],Id_Pc_Add4[21],Id_Pc_Add4[20],
                      Id_Pc_Add4[19],Id_Pc_Add4[18],Id_Pc_Add4[17],
                      Id_Pc_Add4[16],Id_Pc_Add4[15],Id_Pc_Add4[14],
                      Id_Pc_Add4[13],Id_Pc_Add4[12],Id_Pc_Add4[11],
                      Id_Pc_Add4[10],Id_Pc_Add4[9],Id_Pc_Add4[8],Id_Pc_Add4[7],
                      Id_Pc_Add4[6],Id_Pc_Add4[5],Id_Pc_Add4[4],Id_Pc_Add4[3],
                      Id_Pc_Add4[2]}), .px3444 (nx59962z2), .p_EN_int (EN_int), 
                      .p_CLK_int (CLK_int), .px2857 (nx57674z45)) ;
    ALU_0 alu (.p_nbus_Wb_Alu_R ({Wb_Alu_R[31],Wb_Alu_R[30],Wb_Alu_R[29],
          Wb_Alu_R[28],Wb_Alu_R[27],Wb_Alu_R[26],Wb_Alu_R[25],Wb_Alu_R[24],
          Wb_Alu_R[23],Wb_Alu_R[22],Wb_Alu_R[21],Wb_Alu_R[20],Wb_Alu_R[19],
          Wb_Alu_R[18],Wb_Alu_R[17],Wb_Alu_R[16],Wb_Alu_R[15],Wb_Alu_R[14],
          Wb_Alu_R[12],Wb_Alu_R[11],Wb_Alu_R[10],Wb_Alu_R[9],Wb_Alu_R[8],
          Wb_Alu_R[7],Wb_Alu_R[6],Wb_Alu_R[1],Wb_Alu_R[5],Wb_Alu_R[4],
          Wb_Alu_R[3],Wb_Alu_R[2],Wb_Alu_R[13],Wb_Alu_R[0]}), .p_nbus_Wb_D ({
          Wb_D[31],Wb_D[30],Wb_D[29],Wb_D[28],Wb_D[27],Wb_D[26],Wb_D[25],
          Wb_D[24],Wb_D[23],Wb_D[22],Wb_D[21],Wb_D[20],Wb_D[19],Wb_D[18],
          Wb_D[17],Wb_D[16],Wb_D[15],Wb_D[14],Wb_D[12],Wb_D[11],Wb_D[10],Wb_D[9]
          ,Wb_D[8],Wb_D[7],Wb_D[6],Wb_D[1],Wb_D[5],Wb_D[4],Wb_D[3],Wb_D[2],
          Wb_D[13],Wb_D[0]}), .p_nbus_Ex_D2 ({Ex_D2[6],Ex_D2[5],Ex_D2[0],
          Ex_D2[7],Ex_D2[8],Ex_D2[9],Ex_D2[10],Ex_D2[13],Ex_D2[14],Ex_D2[15],
          Ex_D2[16],Ex_D2[17],Ex_D2[18],Ex_D2[19],Ex_D2[20],Ex_D2[21],Ex_D2[22],
          Ex_D2[23],Ex_D2[24],Ex_D2[25],Ex_D2[26],Ex_D2[27],Ex_D2[28],Ex_D2[29],
          Ex_D2[30],Ex_D2[31]}), .\p_Ex_Op(0)   (\Ex_Op(0)  ), .px3439 (
          nx23941z12), .px3432 (nx23941z11), .px3428 (nx23941z10), .px3424 (
          nx23941z9), .px3420 (nx23941z8), .p_nbus_Ex_D1 ({Ex_D1[0],Ex_D1[1],
          Ex_D1[2],Ex_D1[3],Ex_D1[4],Ex_D1[5],Ex_D1[6],Ex_D1[7],Ex_D1[8],
          Ex_D1[9],Ex_D1[10],Ex_D1[11],Ex_D1[12],Ex_D1[13],Ex_D1[14],Ex_D1[15],
          Ex_D1[16],Ex_D1[17],Ex_D1[18],Ex_D1[19],Ex_D1[20],Ex_D1[21],Ex_D1[22],
          Ex_D1[23],Ex_D1[24],Ex_D1[25],Ex_D1[26],Ex_D1[27],Ex_D1[28],Ex_D1[29],
          Ex_D1[30],Ex_D1[31]}), .p_nbus_Ex_Aluc ({Ex_Aluc[0],Ex_Aluc[1],
          Ex_Aluc[2]}), .p_nbus_Mem_Alu_R ({Mem_Alu_R[0],Mem_Alu_R[1],
          Mem_Alu_R[2],Mem_Alu_R[3],Mem_Alu_R[4],Mem_Alu_R[5],Mem_Alu_R[6],
          Mem_Alu_R[7],Mem_Alu_R[8],Mem_Alu_R[9],Mem_Alu_R[10],Mem_Alu_R[11],
          Mem_Alu_R[12],Mem_Alu_R[13],Mem_Alu_R[14],Mem_Alu_R[15],Mem_Alu_R[16],
          Mem_Alu_R[17],Mem_Alu_R[18],Mem_Alu_R[19],Mem_Alu_R[20],Mem_Alu_R[21],
          Mem_Alu_R[22],Mem_Alu_R[23],Mem_Alu_R[24],Mem_Alu_R[25],Mem_Alu_R[26],
          Mem_Alu_R[27],Mem_Alu_R[28],Mem_Alu_R[29],Mem_Alu_R[30],Mem_Alu_R[31]}
          ), .\p_Ex_Extimm(13)   (\Ex_Extimm(13)  ), .px3343 (nx23941z16), .p_nbus_Ex_Fwd_B (
          {Ex_Fwd_B[0],Ex_Fwd_B[1]}), .px3041 (nx30553z1), .px3430 (nx23941z5), 
          .px3040 (nx29556z1), .px3426 (nx23941z4), .px3039 (nx28559z1), .px3422 (
          nx23941z3), .px3038 (nx27562z1), .px3037 (nx26565z1), .px3368 (
          nx57674z1), .px3369 (nx57674z2), .px3030 (nx54097z51), .px3365 (
          nx57674z3), .px3029 (nx54097z52), .px3362 (nx57674z4), .px3028 (
          nx54097z53), .px3359 (nx57674z5), .px3027 (nx54097z54), .px3356 (
          nx57674z6), .px3026 (nx54097z55), .px3353 (nx57674z7), .px3025 (
          nx54097z56), .px3349 (nx57674z8), .px3024 (nx54097z57), .px3345 (
          nx57674z9), .px3023 (nx54097z58), .px3341 (nx57674z10), .px3022 (
          nx54097z59), .px3338 (nx57674z11), .px3021 (nx54097z60), .px3335 (
          nx57674z12), .px3020 (nx54097z61), .px3332 (nx57674z13), .px3019 (
          nx54097z62), .px3329 (nx57674z14), .px3018 (nx54097z63), .px3326 (
          nx57674z15), .px3017 (nx54097z64), .px3323 (nx57674z16), .px3016 (
          nx54097z65), .px3320 (nx57674z17), .px3015 (nx54097z66), .px3317 (
          nx57674z18), .px3014 (nx54097z67), .px3314 (nx57674z19), .px3013 (
          nx54097z68), .px3311 (nx57674z20), .px3012 (nx54097z69), .px3308 (
          nx57674z21), .px3011 (nx54097z70), .px3305 (nx57674z22), .px3010 (
          nx54097z71), .px3302 (nx57674z23), .px3009 (nx54097z72), .px3299 (
          nx57674z24), .px3008 (nx54097z73), .px3296 (nx57674z25), .px3007 (
          nx54097z74), .px3293 (nx57674z26), .px3006 (nx54097z75), .px3290 (
          nx57674z27), .px3005 (nx54097z76), .px3435 (nx57674z28), .px3436 (
          nx57674z29), .px3287 (nx57674z30), .px3004 (nx54097z77), .p_Wb_Reg2reg (
          Wb_Reg2reg), .p_Ex_Aluqb (Ex_Aluqb), .\p_Ex_Extimm(0)   (
          \Ex_Extimm(0)  ), .px3370 (nx23941z1), .px3371 (nx23941z2), .px3373 (
          nx54097z1), .px3366 (nx57674z31), .px3457 (nx54097z2), .px3419 (
          nx57674z32), .px3423 (nx57674z33), .px3427 (nx57674z34), .px3431 (
          nx23941z6), .px3462 (nx23941z13), .px3363 (nx54097z38), .px3463 (
          nx54097z3), .px3360 (nx54097z37), .px3464 (nx54097z4), .px3357 (
          nx54097z41), .px3465 (nx54097z5), .px3354 (nx54097z40), .px3466 (
          nx54097z6), .px3350 (nx57674z35), .px3467 (nx54097z7), .px3346 (
          nx57674z36), .px3468 (nx54097z8), .px3469 (nx54097z9), .px3339 (
          nx54097z44), .px3470 (nx54097z10), .px3336 (nx54097z47), .px3471 (
          nx54097z11), .px3333 (nx54097z32), .px3472 (nx54097z12), .px3330 (
          nx54097z39), .px3473 (nx54097z13), .px3327 (nx54097z50), .px3474 (
          nx54097z14), .px3324 (nx54097z43), .px3475 (nx54097z15), .px3321 (
          nx54097z46), .px3476 (nx54097z16), .px3318 (nx54097z45), .px3477 (
          nx54097z17), .px3315 (nx54097z49), .px3478 (nx54097z18), .px3312 (
          nx21854z1), .px3479 (nx54097z19), .px3309 (nx54097z48), .px3480 (
          nx54097z20), .px3306 (nx54097z42), .px3481 (nx54097z21), .px3303 (
          nx54097z36), .px3482 (nx54097z22), .px3300 (nx54097z35), .px3483 (
          nx54097z23), .px3297 (nx54097z34), .px3484 (nx54097z24), .px3294 (
          nx54097z33), .px3485 (nx54097z25), .px3291 (nx54097z31), .px3486 (
          nx54097z26), .px3288 (nx54097z30), .px3487 (nx54097z27), .p_nbus_Ex_Fwd_A (
          {Ex_Fwd_A[0],Ex_Fwd_A[1]}), .px2963 (nx10566z1), .p_Ex_Z (Ex_Z), .px3206 (
          nx57674z37), .px3209 (nx57674z38), .px3210 (nx57674z39), .px3211 (
          nx57674z40), .px3212 (nx57674z41), .px3213 (nx57674z42), .px3214 (
          nx57674z43), .px3215 (nx57674z44), .px2855 (nx15902z32), .px2964 (
          nx11563z1), .px2965 (nx13559z1), .px2966 (nx14556z1), .px2967 (
          nx15553z1), .px2968 (nx16550z1), .px2969 (nx17547z1), .px2970 (
          nx18544z1), .px2971 (nx19541z1), .px2972 (nx20538z1), .px2973 (
          nx21535z1), .px2974 (nx22532z1), .px2975 (nx24528z1), .px2976 (
          nx25525z1), .px2977 (nx26522z1), .px2978 (nx27519z1), .px2979 (
          nx28516z1), .px2980 (nx29513z1), .px2981 (nx30510z1), .px2982 (
          nx31507z1), .px2983 (nx32504z1), .px2984 (nx33501z1), .px2985 (
          nx13165z1), .px2986 (nx14162z1), .px2987 (nx15159z1), .px2988 (
          nx16156z1), .px2989 (nx17153z1), .px2990 (nx18150z1), .px2991 (
          nx19147z1), .px2992 (nx20144z1), .px2993 (nx21141z1), .px2994 (
          nx22138z1), .px2857 (nx57674z45)) ;
    EX_MEM_unfolded0_0 ex_mem (.px3436 (nx57674z29), .p_nbus_Ex_Aluc ({
                       Ex_Aluc[1],Ex_Aluc[2],Ex_Aluc[0]}), .px3435 (nx57674z28)
                       , .p_CLR_N_int (CLR_N_int), .px3373 (nx54097z1), .p_nbus_Ex_D1 (
                       {Ex_D1[0],Ex_D1[1],Ex_D1[7],Ex_D1[8],Ex_D1[9],Ex_D1[10],
                       Ex_D1[11],Ex_D1[12],Ex_D1[13],Ex_D1[14],Ex_D1[15],
                       Ex_D1[16],Ex_D1[17],Ex_D1[18],Ex_D1[19],Ex_D1[20],
                       Ex_D1[21],Ex_D1[22],Ex_D1[23],Ex_D1[24],Ex_D1[25],
                       Ex_D1[26],Ex_D1[27],Ex_D1[28],Ex_D1[29],Ex_D1[30],
                       Ex_D1[31]}), .px3368 (nx57674z1), .p_nbus_Wb_Alu_R ({
                       Wb_Alu_R[1],Wb_Alu_R[11],Wb_Alu_R[12]}), .p_nbus_Wb_D ({
                       Wb_D[1],Wb_D[11],Wb_D[12]}), .px3367 (nx23941z7), .px3457 (
                       nx54097z2), .px3365 (nx57674z3), .px3463 (nx54097z3), .px3464 (
                       nx54097z4), .px3465 (nx54097z5), .px3466 (nx54097z6), .px3351 (
                       nx23941z14), .px3467 (nx54097z7), .px3349 (nx57674z8), .p_nbus_Ex_Fwd_B (
                       {Ex_Fwd_B[0],Ex_Fwd_B[1]}), .p_Wb_Reg2reg (Wb_Reg2reg), .px3347 (
                       nx23941z15), .px3468 (nx54097z8), .px3345 (nx57674z9), .px3469 (
                       nx54097z9), .px3341 (nx57674z10), .px3470 (nx54097z10), .px3471 (
                       nx54097z11), .px3472 (nx54097z12), .px3473 (nx54097z13), 
                       .px3474 (nx54097z14), .px3475 (nx54097z15), .px3476 (
                       nx54097z16), .px3477 (nx54097z17), .px3478 (nx54097z18), 
                       .px3479 (nx54097z19), .px3311 (nx57674z20), .px3480 (
                       nx54097z20), .px3481 (nx54097z21), .px3482 (nx54097z22), 
                       .px3483 (nx54097z23), .px3484 (nx54097z24), .px3485 (
                       nx54097z25), .px3486 (nx54097z26), .p_nbus_Ex_Fwd_A ({
                       Ex_Fwd_A[0],Ex_Fwd_A[1]}), .px3487 (nx54097z27), .\p_Rt_1_0(0)   (
                       \Rt_1_0(0)  ), .\p_Rt_1_0(1)   (\Rt_1_0(1)  ), .\p_Rt_1_0(2)   (
                       \Rt_1_0(2)  ), .px3258 (nx54097z28), .px3256 (nx23941z18)
                       , .\p_Rs_1_0(1)   (\Rs_1_0(1)  ), .\p_Rs_1_0(0)   (
                       \Rs_1_0(0)  ), .\p_Rs_1_0(2)   (\Rs_1_0(2)  ), .px3255 (
                       nx54097z29), .px3253 (nx23941z17), .px3287 (nx57674z30), 
                       .px3288 (nx54097z30), .px3290 (nx57674z27), .px3291 (
                       nx54097z31), .px3332 (nx57674z13), .px3333 (nx54097z32), 
                       .px3215 (nx57674z44), .px3293 (nx57674z26), .px3294 (
                       nx54097z33), .px3296 (nx57674z25), .px3297 (nx54097z34), 
                       .px3299 (nx57674z24), .px3300 (nx54097z35), .px3214 (
                       nx57674z43), .px3302 (nx57674z23), .px3303 (nx54097z36), 
                       .px3359 (nx57674z5), .px3360 (nx54097z37), .px3362 (
                       nx57674z4), .px3363 (nx54097z38), .px3213 (nx57674z42), .px3329 (
                       nx57674z14), .px3330 (nx54097z39), .px3353 (nx57674z7), .px3354 (
                       nx54097z40), .px3356 (nx57674z6), .px3357 (nx54097z41), .px3212 (
                       nx57674z41), .px3305 (nx57674z22), .px3306 (nx54097z42), 
                       .px3323 (nx57674z16), .px3324 (nx54097z43), .px3338 (
                       nx57674z11), .px3339 (nx54097z44), .px3211 (nx57674z40), 
                       .px3317 (nx57674z18), .px3318 (nx54097z45), .px3320 (
                       nx57674z17), .px3321 (nx54097z46), .px3335 (nx57674z12), 
                       .px3336 (nx54097z47), .px3210 (nx57674z39), .px3308 (
                       nx57674z21), .px3309 (nx54097z48), .px3314 (nx57674z19), 
                       .px3315 (nx54097z49), .px3326 (nx57674z15), .px3327 (
                       nx54097z50), .px3209 (nx57674z38), .p_Ex_Wreg (Ex_Wreg), 
                       .p_Mem_Wreg (Mem_Wreg), .p_Ex_Reg2reg (Ex_Reg2reg), .p_Mem_Reg2reg (
                       Mem_Reg2reg), .p_Ex_Wmem (Ex_Wmem), .p_Mem_Wmem (Mem_Wmem
                       ), .p_nbus_Ex_Rd ({Ex_Rd[0],Ex_Rd[1],Ex_Rd[2]}), .p_nbus_Mem_Rd (
                       {Mem_Rd[0],Mem_Rd[1],Mem_Rd[2]}), .px3030 (nx54097z51), .p_nbus_Mem_Alu_R (
                       {Mem_Alu_R[0],Mem_Alu_R[1],Mem_Alu_R[7],Mem_Alu_R[8],
                       Mem_Alu_R[9],Mem_Alu_R[10],Mem_Alu_R[11],Mem_Alu_R[12],
                       Mem_Alu_R[13],Mem_Alu_R[14],Mem_Alu_R[15],Mem_Alu_R[16],
                       Mem_Alu_R[17],Mem_Alu_R[18],Mem_Alu_R[19],Mem_Alu_R[20],
                       Mem_Alu_R[21],Mem_Alu_R[22],Mem_Alu_R[23],Mem_Alu_R[24],
                       Mem_Alu_R[25],Mem_Alu_R[26],Mem_Alu_R[27],Mem_Alu_R[28],
                       Mem_Alu_R[29],Mem_Alu_R[30],Mem_Alu_R[31]}), .px3029 (
                       nx54097z52), .px3028 (nx54097z53), .px3027 (nx54097z54), 
                       .px3026 (nx54097z55), .px3025 (nx54097z56), .px3024 (
                       nx54097z57), .px3023 (nx54097z58), .px3022 (nx54097z59), 
                       .px3021 (nx54097z60), .px3020 (nx54097z61), .px3019 (
                       nx54097z62), .px3018 (nx54097z63), .px3017 (nx54097z64), 
                       .px3016 (nx54097z65), .px3015 (nx54097z66), .px3014 (
                       nx54097z67), .px3013 (nx54097z68), .px3012 (nx54097z69), 
                       .px3011 (nx54097z70), .px3010 (nx54097z71), .px3009 (
                       nx54097z72), .px3008 (nx54097z73), .px3007 (nx54097z74), 
                       .px3006 (nx54097z75), .px3005 (nx54097z76), .px3004 (
                       nx54097z77), .p_nbus_Ex_D2 ({Ex_D2[0],Ex_D2[1],Ex_D2[2],
                       Ex_D2[3],Ex_D2[4],Ex_D2[5],Ex_D2[6],Ex_D2[7],Ex_D2[8],
                       Ex_D2[9],Ex_D2[10],Ex_D2[11],Ex_D2[12],Ex_D2[13],
                       Ex_D2[14],Ex_D2[15],Ex_D2[16],Ex_D2[17],Ex_D2[18],
                       Ex_D2[19],Ex_D2[20],Ex_D2[21],Ex_D2[22],Ex_D2[23],
                       Ex_D2[24],Ex_D2[25],Ex_D2[26],Ex_D2[27],Ex_D2[28],
                       Ex_D2[29],Ex_D2[30],Ex_D2[31]}), .p_nbus_Mem_D2 ({
                       Mem_D2[0],Mem_D2[1],Mem_D2[2],Mem_D2[3],Mem_D2[4],
                       Mem_D2[5],Mem_D2[6],Mem_D2[7],Mem_D2[8],Mem_D2[9],
                       Mem_D2[10],Mem_D2[11],Mem_D2[12],Mem_D2[13],Mem_D2[14],
                       Mem_D2[15],Mem_D2[16],Mem_D2[17],Mem_D2[18],Mem_D2[19],
                       Mem_D2[20],Mem_D2[21],Mem_D2[22],Mem_D2[23],Mem_D2[24],
                       Mem_D2[25],Mem_D2[26],Mem_D2[27],Mem_D2[28],Mem_D2[29],
                       Mem_D2[30],Mem_D2[31]}), .px3433 (nx58593z1), .p_EN_int (
                       EN_int), .p_CLK_int (CLK_int)) ;
    DATAMEM_unfolded0_0 data_mem (.p_rtlcs428 (nx22656z1), .px3406 (nx4630z1), .p_rtlcs427 (
                        nx22656z2), .px3405 (nx3633z1), .p_rtlcs426 (nx22656z3)
                        , .px3404 (nx1637z1), .p_rtlcs425 (nx22656z4), .px3403 (
                        nx640z1), .p_rtlcs424 (nx22656z5), .px3402 (nx65179z1), 
                        .p_rtlcs423 (nx22656z6), .px3401 (nx64182z1), .p_rtlcs422 (
                        nx22656z7), .px3400 (nx63185z1), .p_rtlcs421 (nx22656z8)
                        , .px3399 (nx62188z1), .p_rtlcs420 (nx22656z9), .px3398 (
                        nx61191z1), .p_rtlcs419 (nx22656z10), .px3397 (nx60194z1
                        ), .p_rtlcs418 (nx22656z11), .px3396 (nx59197z1), .p_rtlcs417 (
                        nx22656z12), .px3395 (nx58200z1), .p_rtlcs416 (
                        nx22656z13), .px3394 (nx56204z1), .p_rtlcs415 (
                        nx22656z14), .px3393 (nx55207z1), .p_rtlcs414 (
                        nx22656z15), .px3392 (nx54210z1), .p_rtlcs413 (
                        nx22656z16), .px3391 (nx53213z1), .p_rtlcs412 (
                        nx22656z17), .px3390 (nx52216z1), .p_rtlcs411 (
                        nx22656z18), .px3389 (nx51219z1), .p_rtlcs410 (
                        nx22656z19), .px3388 (nx50222z1), .p_rtlcs409 (
                        nx22656z20), .px3387 (nx49225z1), .p_rtlcs408 (
                        nx22656z21), .px3386 (nx48228z1), .p_rtlcs407 (
                        nx22656z22), .px3385 (nx47231z1), .p_rtlcs406 (
                        nx22656z23), .px3384 (nx7359z1), .p_rtlcs405 (nx22656z24
                        ), .px3383 (nx6362z1), .p_rtlcs404 (nx22656z25), .px3382 (
                        nx5365z1), .p_rtlcs403 (nx22656z26), .px3381 (nx4368z1)
                        , .p_rtlcs402 (nx22656z27), .px3380 (nx3371z1), .p_rtlcs401 (
                        nx22656z28), .px3379 (nx2374z1), .p_rtlcs400 (nx22656z29
                        ), .px3378 (nx1377z1), .p_rtlcs399 (nx22656z30), .px3377 (
                        nx380z1), .p_rtlcs398 (nx22656z31), .px3376 (nx64919z1)
                        , .p_rtlcs397 (nx22656z32), .px3375 (nx63922z1), .px3455 (
                        nx60794z1), .p_nbus_Mem_Alu_R ({Mem_Alu_R[2],
                        Mem_Alu_R[3],Mem_Alu_R[4],Mem_Alu_R[5],Mem_Alu_R[6]}), .p_CLR_N_int (
                        CLR_N_int), .p_pc_not_clr_n (pc_not_clr_n), .p_Mem_Wmem (
                        Mem_Wmem), .p_CLK_int (CLK_int)) ;
    BUFGP CLK_ibuf (.O (CLK_int), .I (CLK)) ;
endmodule


module DATAMEM_unfolded0_0 ( p_rtlcs428, px3406, p_rtlcs427, px3405, p_rtlcs426, 
                             px3404, p_rtlcs425, px3403, p_rtlcs424, px3402, 
                             p_rtlcs423, px3401, p_rtlcs422, px3400, p_rtlcs421, 
                             px3399, p_rtlcs420, px3398, p_rtlcs419, px3397, 
                             p_rtlcs418, px3396, p_rtlcs417, px3395, p_rtlcs416, 
                             px3394, p_rtlcs415, px3393, p_rtlcs414, px3392, 
                             p_rtlcs413, px3391, p_rtlcs412, px3390, p_rtlcs411, 
                             px3389, p_rtlcs410, px3388, p_rtlcs409, px3387, 
                             p_rtlcs408, px3386, p_rtlcs407, px3385, p_rtlcs406, 
                             px3384, p_rtlcs405, px3383, p_rtlcs404, px3382, 
                             p_rtlcs403, px3381, p_rtlcs402, px3380, p_rtlcs401, 
                             px3379, p_rtlcs400, px3378, p_rtlcs399, px3377, 
                             p_rtlcs398, px3376, p_rtlcs397, px3375, px3455, 
                             p_nbus_Mem_Alu_R, p_CLR_N_int, p_pc_not_clr_n, 
                             p_Mem_Wmem, p_CLK_int ) ;

    input p_rtlcs428 ;
    output px3406 ;
    input p_rtlcs427 ;
    output px3405 ;
    input p_rtlcs426 ;
    output px3404 ;
    input p_rtlcs425 ;
    output px3403 ;
    input p_rtlcs424 ;
    output px3402 ;
    input p_rtlcs423 ;
    output px3401 ;
    input p_rtlcs422 ;
    output px3400 ;
    input p_rtlcs421 ;
    output px3399 ;
    input p_rtlcs420 ;
    output px3398 ;
    input p_rtlcs419 ;
    output px3397 ;
    input p_rtlcs418 ;
    output px3396 ;
    input p_rtlcs417 ;
    output px3395 ;
    input p_rtlcs416 ;
    output px3394 ;
    input p_rtlcs415 ;
    output px3393 ;
    input p_rtlcs414 ;
    output px3392 ;
    input p_rtlcs413 ;
    output px3391 ;
    input p_rtlcs412 ;
    output px3390 ;
    input p_rtlcs411 ;
    output px3389 ;
    input p_rtlcs410 ;
    output px3388 ;
    input p_rtlcs409 ;
    output px3387 ;
    input p_rtlcs408 ;
    output px3386 ;
    input p_rtlcs407 ;
    output px3385 ;
    input p_rtlcs406 ;
    output px3384 ;
    input p_rtlcs405 ;
    output px3383 ;
    input p_rtlcs404 ;
    output px3382 ;
    input p_rtlcs403 ;
    output px3381 ;
    input p_rtlcs402 ;
    output px3380 ;
    input p_rtlcs401 ;
    output px3379 ;
    input p_rtlcs400 ;
    output px3378 ;
    input p_rtlcs399 ;
    output px3377 ;
    input p_rtlcs398 ;
    output px3376 ;
    input p_rtlcs397 ;
    output px3375 ;
    output px3455 ;
    input [31:27]p_nbus_Mem_Alu_R ;
    input p_CLR_N_int ;
    output p_pc_not_clr_n ;
    input p_Mem_Wmem ;
    input p_CLK_int ;

    wire nx11305z6, nx11305z5, nx11305z4, nx11305z3, nx11305z11, nx11305z10, 
         nx11305z9, nx11305z8, nx11305z7, nx11305z2, nx39150z1;
    wire [0:31]data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3;
    wire nx38153z1, nx37156z1, nx36159z1, nx35162z1, nx34165z1, nx33168z1, 
         nx32171z1, nx31174z1, nx30177z1, nx20641z1, nx19644z1, nx18647z1, 
         nx17650z1, nx16653z1, nx15656z1, nx14659z1, nx13662z1, nx12665z1, 
         nx11668z1, nx9672z1, nx8675z1, nx7678z1, nx6681z1, nx5684z1, nx4687z1, 
         nx3690z1, nx2693z1, nx1696z1, nx699z1, nx64239z1, nx63242z1, nx6, nx7, 
         nx45, nx47, nx49, nx51, nx53, nx55, nx57, nx59, nx61, nx63, nx65, nx67, 
         nx69, nx71, nx73, nx75, nx77, nx79, nx81, nx83, nx85, nx87, nx89, nx91, 
         nx93, nx95, nx97, nx99, nx101, nx103, nx105;



    INV ix9672z1317 (.O (p_pc_not_clr_n), .I (p_CLR_N_int)) ;
    LUT6 ix39150z1314 (.O (nx39150z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix39150z1314.INIT = 64'h0000000100000000;
    LUT6 ix38153z1314 (.O (nx38153z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix38153z1314.INIT = 64'h0001000000000000;
    LUT6 ix37156z1314 (.O (nx37156z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix37156z1314.INIT = 64'h0000010000000000;
    LUT6 ix36159z1314 (.O (nx36159z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix36159z1314.INIT = 64'h0100000000000000;
    LUT6 ix35162z1314 (.O (nx35162z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix35162z1314.INIT = 64'h0000001000000000;
    LUT6 ix34165z1314 (.O (nx34165z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix34165z1314.INIT = 64'h0010000000000000;
    LUT6 ix33168z1314 (.O (nx33168z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix33168z1314.INIT = 64'h0000100000000000;
    LUT6 ix32171z1314 (.O (nx32171z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix32171z1314.INIT = 64'h1000000000000000;
    LUT6 ix31174z1314 (.O (nx31174z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix31174z1314.INIT = 64'h0000000400000000;
    LUT6 ix30177z1314 (.O (nx30177z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix30177z1314.INIT = 64'h0004000000000000;
    LUT6 ix20641z1314 (.O (nx20641z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix20641z1314.INIT = 64'h0000040000000000;
    LUT6 ix19644z1314 (.O (nx19644z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix19644z1314.INIT = 64'h0400000000000000;
    LUT6 ix18647z1314 (.O (nx18647z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix18647z1314.INIT = 64'h0000004000000000;
    LUT6 ix17650z1314 (.O (nx17650z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix17650z1314.INIT = 64'h0040000000000000;
    LUT6 ix16653z1314 (.O (nx16653z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix16653z1314.INIT = 64'h0000400000000000;
    LUT6 ix15656z1314 (.O (nx15656z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix15656z1314.INIT = 64'h4000000000000000;
    LUT6 ix14659z1314 (.O (nx14659z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix14659z1314.INIT = 64'h0000000200000000;
    LUT6 ix13662z1314 (.O (nx13662z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix13662z1314.INIT = 64'h0002000000000000;
    LUT6 ix12665z1314 (.O (nx12665z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix12665z1314.INIT = 64'h0000020000000000;
    LUT6 ix11668z1314 (.O (nx11668z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix11668z1314.INIT = 64'h0200000000000000;
    LUT6 ix9672z1314 (.O (nx9672z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix9672z1314.INIT = 64'h0000002000000000;
    LUT6 ix8675z1314 (.O (nx8675z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix8675z1314.INIT = 64'h0020000000000000;
    LUT6 ix7678z1314 (.O (nx7678z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix7678z1314.INIT = 64'h0000200000000000;
    LUT6 ix6681z1314 (.O (nx6681z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix6681z1314.INIT = 64'h2000000000000000;
    LUT6 ix5684z1314 (.O (nx5684z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix5684z1314.INIT = 64'h0000000800000000;
    LUT6 ix4687z1314 (.O (nx4687z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix4687z1314.INIT = 64'h0008000000000000;
    LUT6 ix3690z1314 (.O (nx3690z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix3690z1314.INIT = 64'h0000080000000000;
    LUT6 ix2693z1314 (.O (nx2693z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix2693z1314.INIT = 64'h0800000000000000;
    LUT6 ix1696z1314 (.O (nx1696z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix1696z1314.INIT = 64'h0000008000000000;
    LUT6 ix699z1314 (.O (nx699z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix699z1314.INIT = 64'h0080000000000000;
    LUT6 ix64239z1314 (.O (nx64239z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix64239z1314.INIT = 64'h0000800000000000;
    LUT6 ix63242z1314 (.O (nx63242z1), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Mem_Alu_R[29]), .I3 (
         p_nbus_Mem_Alu_R[30]), .I4 (p_nbus_Mem_Alu_R[31]), .I5 (px3455)) ;
         defparam ix63242z1314.INIT = 64'h8000000000000000;
    (* HLUTNM = "LUT62_6_4" *)
    LUT4 ix7314z45346 (.O (px3375), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs397)) ;
         defparam ix7314z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_5" *)
    LUT4 ix7315z45346 (.O (px3376), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs398)) ;
         defparam ix7315z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_5" *)
    LUT4 ix7316z45346 (.O (px3377), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs399)) ;
         defparam ix7316z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_6" *)
    LUT4 ix7317z45346 (.O (px3378), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs400)) ;
         defparam ix7317z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_6" *)
    LUT4 ix7318z45346 (.O (px3379), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs401)) ;
         defparam ix7318z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_7" *)
    LUT4 ix8306z45346 (.O (px3380), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs402)) ;
         defparam ix8306z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_7" *)
    LUT4 ix8307z45346 (.O (px3381), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs403)) ;
         defparam ix8307z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_8" *)
    LUT4 ix8308z45346 (.O (px3382), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs404)) ;
         defparam ix8308z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_8" *)
    LUT4 ix8309z45346 (.O (px3383), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs405)) ;
         defparam ix8309z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_9" *)
    LUT4 ix8310z45346 (.O (px3384), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs406)) ;
         defparam ix8310z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_9" *)
    LUT4 ix8311z45346 (.O (px3385), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs407)) ;
         defparam ix8311z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_10" *)
    LUT4 ix8312z45346 (.O (px3386), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs408)) ;
         defparam ix8312z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_10" *)
    LUT4 ix8313z45346 (.O (px3387), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs409)) ;
         defparam ix8313z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_11" *)
    LUT4 ix8314z45346 (.O (px3388), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs410)) ;
         defparam ix8314z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_11" *)
    LUT4 ix8315z45346 (.O (px3389), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs411)) ;
         defparam ix8315z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_12" *)
    LUT4 ix9303z45346 (.O (px3390), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs412)) ;
         defparam ix9303z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_12" *)
    LUT4 ix9304z45346 (.O (px3391), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs413)) ;
         defparam ix9304z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_13" *)
    LUT4 ix9305z45346 (.O (px3392), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs414)) ;
         defparam ix9305z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_13" *)
    LUT4 ix9306z45346 (.O (px3393), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs415)) ;
         defparam ix9306z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_14" *)
    LUT4 ix9307z45346 (.O (px3394), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs416)) ;
         defparam ix9307z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_14" *)
    LUT4 ix9308z45346 (.O (px3395), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs417)) ;
         defparam ix9308z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_15" *)
    LUT4 ix9309z45346 (.O (px3396), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs418)) ;
         defparam ix9309z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_15" *)
    LUT4 ix9310z45346 (.O (px3397), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs419)) ;
         defparam ix9310z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_16" *)
    LUT4 ix9311z45346 (.O (px3398), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs420)) ;
         defparam ix9311z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_16" *)
    LUT4 ix9312z45346 (.O (px3399), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs421)) ;
         defparam ix9312z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_1" *)
    LUT4 ix11299z45346 (.O (px3400), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs422)) ;
         defparam ix11299z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_1" *)
    LUT4 ix11300z45346 (.O (px3401), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs423)) ;
         defparam ix11300z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_2" *)
    LUT4 ix11301z45346 (.O (px3402), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs424)) ;
         defparam ix11301z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_2" *)
    LUT4 ix11302z45346 (.O (px3403), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs425)) ;
         defparam ix11302z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_3" *)
    LUT4 ix11303z45346 (.O (px3404), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs426)) ;
         defparam ix11303z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_3" *)
    LUT4 ix11304z45346 (.O (px3405), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs427)) ;
         defparam ix11304z45346.INIT = 16'hAC00;
    (* HLUTNM = "LUT62_6_4" *)
    LUT4 ix11305z45346 (.O (px3406), .I0 (nx11305z2), .I1 (nx11305z7), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_rtlcs428)) ;
         defparam ix11305z45346.INIT = 16'hAC00;
    LUT6 ix11305z53748 (.O (nx11305z7), .I0 (nx11305z8), .I1 (nx11305z9), .I2 (
         nx11305z10), .I3 (nx11305z11), .I4 (p_nbus_Mem_Alu_R[28]), .I5 (
         p_nbus_Mem_Alu_R[29])) ;
         defparam ix11305z53748.INIT = 64'hF0F0AAAAFF00CCCC;
    LUT6 ix11305z45339 (.O (nx11305z11), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[8]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[9]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[10]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[11])) ;
         defparam ix11305z45339.INIT = 64'h0145236789CDABEF;
    LUT6 ix11305z45338 (.O (nx11305z10), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[12]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[13]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[14]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[15])) ;
         defparam ix11305z45338.INIT = 64'h0145236789CDABEF;
    LUT6 ix11305z45337 (.O (nx11305z9), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[0]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[1]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[2]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[3])) ;
         defparam ix11305z45337.INIT = 64'h0145236789CDABEF;
    LUT6 ix11305z45336 (.O (nx11305z8), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[4]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[5]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[6]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[7])) ;
         defparam ix11305z45336.INIT = 64'h0145236789CDABEF;
    LUT6 ix11305z53743 (.O (nx11305z2), .I0 (nx11305z3), .I1 (nx11305z4), .I2 (
         nx11305z5), .I3 (nx11305z6), .I4 (p_nbus_Mem_Alu_R[28]), .I5 (
         p_nbus_Mem_Alu_R[29])) ;
         defparam ix11305z53743.INIT = 64'hF0F0AAAAFF00CCCC;
    LUT6 ix11305z45334 (.O (nx11305z6), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[24]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[25]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[26]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[27])) ;
         defparam ix11305z45334.INIT = 64'h0145236789CDABEF;
    LUT6 ix11305z45333 (.O (nx11305z5), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[28]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[29]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[30]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[31])) ;
         defparam ix11305z45333.INIT = 64'h0145236789CDABEF;
    LUT6 ix11305z45332 (.O (nx11305z4), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[16]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[17]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[18]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[19])) ;
         defparam ix11305z45332.INIT = 64'h0145236789CDABEF;
    LUT6 ix11305z45331 (.O (nx11305z3), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[20]), .I3 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[21]), .I4 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[22]), .I5 (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[23])) ;
         defparam ix11305z45331.INIT = 64'h0145236789CDABEF;
    LUT2 ix9672z1323 (.O (px3455), .I0 (p_Mem_Wmem), .I1 (p_CLR_N_int)) ;
         defparam ix9672z1323.INIT = 4'h8;
    VCC \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(31)_I21_FD_PWR  (.P (
        nx6)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(31)_I21_FD_LUT  (.O (
         nx7), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[31]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[31]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(31)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(31)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[31]), .C (
         p_CLK_int), .CE (nx6), .D (nx7), .R (nx63242z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(30)_I21_FD_LUT  (.O (
         nx45), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[30])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[30]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(30)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(30)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[30]), .C (
         p_CLK_int), .CE (nx6), .D (nx45), .R (nx64239z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(29)_I21_FD_LUT  (.O (
         nx47), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[29])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[29]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(29)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(29)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[29]), .C (
         p_CLK_int), .CE (nx6), .D (nx47), .R (nx699z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(28)_I21_FD_LUT  (.O (
         nx49), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[28])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[28]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(28)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(28)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[28]), .C (
         p_CLK_int), .CE (nx6), .D (nx49), .R (nx1696z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(27)_I21_FD_LUT  (.O (
         nx51), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[27])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[27]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(27)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(27)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[27]), .C (
         p_CLK_int), .CE (nx6), .D (nx51), .R (nx2693z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(26)_I21_FD_LUT  (.O (
         nx53), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[26])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[26]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(26)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(26)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[26]), .C (
         p_CLK_int), .CE (nx6), .D (nx53), .R (nx3690z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(25)_I21_FD_LUT  (.O (
         nx55), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[25])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[25]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(25)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(25)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[25]), .C (
         p_CLK_int), .CE (nx6), .D (nx55), .R (nx4687z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(24)_I21_FD_LUT  (.O (
         nx57), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[24])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[24]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(24)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(24)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[24]), .C (
         p_CLK_int), .CE (nx6), .D (nx57), .R (nx5684z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(23)_I21_FD_LUT  (.O (
         nx59), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[23])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[23]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(23)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(23)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[23]), .C (
         p_CLK_int), .CE (nx6), .D (nx59), .R (nx6681z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(22)_I21_FD_LUT  (.O (
         nx61), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[22])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[22]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(22)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(22)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[22]), .C (
         p_CLK_int), .CE (nx6), .D (nx61), .R (nx7678z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(21)_I21_FD_LUT  (.O (
         nx63), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[21])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[21]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(21)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(21)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[21]), .C (
         p_CLK_int), .CE (nx6), .D (nx63), .R (nx8675z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(20)_I21_FD_LUT  (.O (
         nx65), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[20])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[20]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(20)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(20)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[20]), .C (
         p_CLK_int), .CE (nx6), .D (nx65), .R (nx9672z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(19)_I21_FD_LUT  (.O (
         nx67), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[19])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[19]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(19)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(19)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[19]), .C (
         p_CLK_int), .CE (nx6), .D (nx67), .R (nx11668z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(18)_I21_FD_LUT  (.O (
         nx69), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[18])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[18]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(18)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(18)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[18]), .C (
         p_CLK_int), .CE (nx6), .D (nx69), .R (nx12665z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(17)_I21_FD_LUT  (.O (
         nx71), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[17])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[17]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(17)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(17)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[17]), .C (
         p_CLK_int), .CE (nx6), .D (nx71), .R (nx13662z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(16)_I21_FD_LUT  (.O (
         nx73), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[16])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[16]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(16)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(16)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[16]), .C (
         p_CLK_int), .CE (nx6), .D (nx73), .R (nx14659z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(15)_I21_FD_LUT  (.O (
         nx75), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[15])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[15]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(15)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(15)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[15]), .C (
         p_CLK_int), .CE (nx6), .D (nx75), .R (nx15656z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(14)_I21_FD_LUT  (.O (
         nx77), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[14])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[14]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(14)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(14)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[14]), .C (
         p_CLK_int), .CE (nx6), .D (nx77), .R (nx16653z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(13)_I21_FD_LUT  (.O (
         nx79), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[13])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[13]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(13)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(13)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[13]), .C (
         p_CLK_int), .CE (nx6), .D (nx79), .R (nx17650z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(12)_I21_FD_LUT  (.O (
         nx81), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[12])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[12]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(12)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(12)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[12]), .C (
         p_CLK_int), .CE (nx6), .D (nx81), .R (nx18647z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(11)_I21_FD_LUT  (.O (
         nx83), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[11])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[11]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(11)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(11)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[11]), .C (
         p_CLK_int), .CE (nx6), .D (nx83), .R (nx19644z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(10)_I21_FD_LUT  (.O (
         nx85), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[10])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[10]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(10)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(10)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[10]), .C (
         p_CLK_int), .CE (nx6), .D (nx85), .R (nx20641z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(9)_I21_FD_LUT  (.O (
         nx87), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[9]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[9]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(9)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(9)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[9]), .C (
         p_CLK_int), .CE (nx6), .D (nx87), .R (nx30177z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(8)_I21_FD_LUT  (.O (
         nx89), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[8]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[8]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(8)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(8)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[8]), .C (
         p_CLK_int), .CE (nx6), .D (nx89), .R (nx31174z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(7)_I21_FD_LUT  (.O (
         nx91), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[7]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[7]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(7)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(7)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[7]), .C (
         p_CLK_int), .CE (nx6), .D (nx91), .R (nx32171z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(6)_I21_FD_LUT  (.O (
         nx93), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[6]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[6]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(6)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(6)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[6]), .C (
         p_CLK_int), .CE (nx6), .D (nx93), .R (nx33168z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(5)_I21_FD_LUT  (.O (
         nx95), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[5]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[5]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(5)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(5)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[5]), .C (
         p_CLK_int), .CE (nx6), .D (nx95), .R (nx34165z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(4)_I21_FD_LUT  (.O (
         nx97), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[4]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[4]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(4)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(4)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[4]), .C (
         p_CLK_int), .CE (nx6), .D (nx97), .R (nx35162z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(3)_I21_FD_LUT  (.O (
         nx99), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[3]), 
         .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[3]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(3)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(3)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[3]), .C (
         p_CLK_int), .CE (nx6), .D (nx99), .R (nx36159z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(2)_I21_FD_LUT  (.O (
         nx101), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[2])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[2]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(2)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(2)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[2]), .C (
         p_CLK_int), .CE (nx6), .D (nx101), .R (nx37156z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(1)_I21_FD_LUT  (.O (
         nx103), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[1])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[1]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(1)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(1)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[1]), .C (
         p_CLK_int), .CE (nx6), .D (nx103), .R (nx38153z1)) ;
    LUT4 \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(0)_I21_FD_LUT  (.O (
         nx105), .I0 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[0])
         , .I1 (data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[0]), .I2 (
         p_Mem_Wmem), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(0)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3(0)  (.Q (
         data_mem_MSR__DATAMEM_ROM_4_rtlc_sync_msr_n0_rtlcGen3[0]), .C (
         p_CLK_int), .CE (nx6), .D (nx105), .R (nx39150z1)) ;
endmodule


module EX_MEM_unfolded0_0 ( px3436, p_nbus_Ex_Aluc, px3435, p_CLR_N_int, px3373, 
                            p_nbus_Ex_D1, px3368, p_nbus_Wb_Alu_R, p_nbus_Wb_D, 
                            px3367, px3457, px3365, px3463, px3464, px3465, 
                            px3466, px3351, px3467, px3349, p_nbus_Ex_Fwd_B, 
                            p_Wb_Reg2reg, px3347, px3468, px3345, px3469, px3341, 
                            px3470, px3471, px3472, px3473, px3474, px3475, 
                            px3476, px3477, px3478, px3479, px3311, px3480, 
                            px3481, px3482, px3483, px3484, px3485, px3486, 
                            p_nbus_Ex_Fwd_A, px3487, \p_Rt_1_0(0)  , 
                            \p_Rt_1_0(1)  , \p_Rt_1_0(2)  , px3258, px3256, 
                            \p_Rs_1_0(1)  , \p_Rs_1_0(0)  , \p_Rs_1_0(2)  , 
                            px3255, px3253, px3287, px3288, px3290, px3291, 
                            px3332, px3333, px3215, px3293, px3294, px3296, 
                            px3297, px3299, px3300, px3214, px3302, px3303, 
                            px3359, px3360, px3362, px3363, px3213, px3329, 
                            px3330, px3353, px3354, px3356, px3357, px3212, 
                            px3305, px3306, px3323, px3324, px3338, px3339, 
                            px3211, px3317, px3318, px3320, px3321, px3335, 
                            px3336, px3210, px3308, px3309, px3314, px3315, 
                            px3326, px3327, px3209, p_Ex_Wreg, p_Mem_Wreg, 
                            p_Ex_Reg2reg, p_Mem_Reg2reg, p_Ex_Wmem, p_Mem_Wmem, 
                            p_nbus_Ex_Rd, p_nbus_Mem_Rd, px3030, 
                            p_nbus_Mem_Alu_R, px3029, px3028, px3027, px3026, 
                            px3025, px3024, px3023, px3022, px3021, px3020, 
                            px3019, px3018, px3017, px3016, px3015, px3014, 
                            px3013, px3012, px3011, px3010, px3009, px3008, 
                            px3007, px3006, px3005, px3004, p_nbus_Ex_D2, 
                            p_nbus_Mem_D2, px3433, p_EN_int, p_CLK_int ) ;

    output px3436 ;
    input [2:0]p_nbus_Ex_Aluc ;
    output px3435 ;
    input p_CLR_N_int ;
    input px3373 ;
    input [31:5]p_nbus_Ex_D1 ;
    output px3368 ;
    input [31:29]p_nbus_Wb_Alu_R ;
    input [31:29]p_nbus_Wb_D ;
    output px3367 ;
    input px3457 ;
    output px3365 ;
    input px3463 ;
    input px3464 ;
    input px3465 ;
    input px3466 ;
    output px3351 ;
    input px3467 ;
    output px3349 ;
    input [1:0]p_nbus_Ex_Fwd_B ;
    input p_Wb_Reg2reg ;
    output px3347 ;
    input px3468 ;
    output px3345 ;
    input px3469 ;
    output px3341 ;
    input px3470 ;
    input px3471 ;
    input px3472 ;
    input px3473 ;
    input px3474 ;
    input px3475 ;
    input px3476 ;
    input px3477 ;
    input px3478 ;
    input px3479 ;
    output px3311 ;
    input px3480 ;
    input px3481 ;
    input px3482 ;
    input px3483 ;
    input px3484 ;
    input px3485 ;
    input px3486 ;
    input [1:0]p_nbus_Ex_Fwd_A ;
    input px3487 ;
    input \p_Rt_1_0(0)   ;
    input \p_Rt_1_0(1)   ;
    input \p_Rt_1_0(2)   ;
    input px3258 ;
    output px3256 ;
    input \p_Rs_1_0(1)   ;
    input \p_Rs_1_0(0)   ;
    input \p_Rs_1_0(2)   ;
    input px3255 ;
    output px3253 ;
    output px3287 ;
    input px3288 ;
    output px3290 ;
    input px3291 ;
    output px3332 ;
    input px3333 ;
    output px3215 ;
    output px3293 ;
    input px3294 ;
    output px3296 ;
    input px3297 ;
    output px3299 ;
    input px3300 ;
    output px3214 ;
    output px3302 ;
    input px3303 ;
    output px3359 ;
    input px3360 ;
    output px3362 ;
    input px3363 ;
    output px3213 ;
    output px3329 ;
    input px3330 ;
    output px3353 ;
    input px3354 ;
    output px3356 ;
    input px3357 ;
    output px3212 ;
    output px3305 ;
    input px3306 ;
    output px3323 ;
    input px3324 ;
    output px3338 ;
    input px3339 ;
    output px3211 ;
    output px3317 ;
    input px3318 ;
    output px3320 ;
    input px3321 ;
    output px3335 ;
    input px3336 ;
    output px3210 ;
    output px3308 ;
    input px3309 ;
    output px3314 ;
    input px3315 ;
    output px3326 ;
    input px3327 ;
    output px3209 ;
    input p_Ex_Wreg ;
    output p_Mem_Wreg ;
    input p_Ex_Reg2reg ;
    output p_Mem_Reg2reg ;
    input p_Ex_Wmem ;
    output p_Mem_Wmem ;
    input [2:0]p_nbus_Ex_Rd ;
    output [2:0]p_nbus_Mem_Rd ;
    input px3030 ;
    output [31:5]p_nbus_Mem_Alu_R ;
    input px3029 ;
    input px3028 ;
    input px3027 ;
    input px3026 ;
    input px3025 ;
    input px3024 ;
    input px3023 ;
    input px3022 ;
    input px3021 ;
    input px3020 ;
    input px3019 ;
    input px3018 ;
    input px3017 ;
    input px3016 ;
    input px3015 ;
    input px3014 ;
    input px3013 ;
    input px3012 ;
    input px3011 ;
    input px3010 ;
    input px3009 ;
    input px3008 ;
    input px3007 ;
    input px3006 ;
    input px3005 ;
    input px3004 ;
    input [31:0]p_nbus_Ex_D2 ;
    output [31:0]p_nbus_Mem_D2 ;
    output px3433 ;
    input p_EN_int ;
    input p_CLK_int ;

    wire nx59888z3, nx59885z3;



    FDRE \reg_Mem_D2(31)  (.Q (p_nbus_Mem_D2[0]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[0]), .R (px3433)) ;
    FDRE \reg_Mem_D2(30)  (.Q (p_nbus_Mem_D2[1]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[1]), .R (px3433)) ;
    FDRE \reg_Mem_D2(29)  (.Q (p_nbus_Mem_D2[2]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[2]), .R (px3433)) ;
    FDRE \reg_Mem_D2(28)  (.Q (p_nbus_Mem_D2[3]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[3]), .R (px3433)) ;
    FDRE \reg_Mem_D2(27)  (.Q (p_nbus_Mem_D2[4]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[4]), .R (px3433)) ;
    FDRE \reg_Mem_D2(26)  (.Q (p_nbus_Mem_D2[5]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[5]), .R (px3433)) ;
    FDRE \reg_Mem_D2(25)  (.Q (p_nbus_Mem_D2[6]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[6]), .R (px3433)) ;
    FDRE \reg_Mem_D2(24)  (.Q (p_nbus_Mem_D2[7]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[7]), .R (px3433)) ;
    FDRE \reg_Mem_D2(23)  (.Q (p_nbus_Mem_D2[8]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[8]), .R (px3433)) ;
    FDRE \reg_Mem_D2(22)  (.Q (p_nbus_Mem_D2[9]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[9]), .R (px3433)) ;
    FDRE \reg_Mem_D2(21)  (.Q (p_nbus_Mem_D2[10]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[10]), .R (px3433)) ;
    FDRE \reg_Mem_D2(20)  (.Q (p_nbus_Mem_D2[11]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[11]), .R (px3433)) ;
    FDRE \reg_Mem_D2(19)  (.Q (p_nbus_Mem_D2[12]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[12]), .R (px3433)) ;
    FDRE \reg_Mem_D2(18)  (.Q (p_nbus_Mem_D2[13]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[13]), .R (px3433)) ;
    FDRE \reg_Mem_D2(17)  (.Q (p_nbus_Mem_D2[14]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[14]), .R (px3433)) ;
    FDRE \reg_Mem_D2(16)  (.Q (p_nbus_Mem_D2[15]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[15]), .R (px3433)) ;
    FDRE \reg_Mem_D2(15)  (.Q (p_nbus_Mem_D2[16]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[16]), .R (px3433)) ;
    FDRE \reg_Mem_D2(14)  (.Q (p_nbus_Mem_D2[17]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[17]), .R (px3433)) ;
    FDRE \reg_Mem_D2(13)  (.Q (p_nbus_Mem_D2[18]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[18]), .R (px3433)) ;
    FDRE \reg_Mem_D2(12)  (.Q (p_nbus_Mem_D2[19]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[19]), .R (px3433)) ;
    FDRE \reg_Mem_D2(11)  (.Q (p_nbus_Mem_D2[20]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[20]), .R (px3433)) ;
    FDRE \reg_Mem_D2(10)  (.Q (p_nbus_Mem_D2[21]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (p_nbus_Ex_D2[21]), .R (px3433)) ;
    FDRE \reg_Mem_D2(9)  (.Q (p_nbus_Mem_D2[22]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[22]), .R (px3433)) ;
    FDRE \reg_Mem_D2(8)  (.Q (p_nbus_Mem_D2[23]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[23]), .R (px3433)) ;
    FDRE \reg_Mem_D2(7)  (.Q (p_nbus_Mem_D2[24]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[24]), .R (px3433)) ;
    FDRE \reg_Mem_D2(6)  (.Q (p_nbus_Mem_D2[25]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[25]), .R (px3433)) ;
    FDRE \reg_Mem_D2(5)  (.Q (p_nbus_Mem_D2[26]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[26]), .R (px3433)) ;
    FDRE \reg_Mem_D2(4)  (.Q (p_nbus_Mem_D2[27]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[27]), .R (px3433)) ;
    FDRE \reg_Mem_D2(3)  (.Q (p_nbus_Mem_D2[28]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[28]), .R (px3433)) ;
    FDRE \reg_Mem_D2(2)  (.Q (p_nbus_Mem_D2[29]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[29]), .R (px3433)) ;
    FDRE \reg_Mem_D2(1)  (.Q (p_nbus_Mem_D2[30]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[30]), .R (px3433)) ;
    FDRE \reg_Mem_D2(0)  (.Q (p_nbus_Mem_D2[31]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_D2[31]), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(31)  (.Q (p_nbus_Mem_Alu_R[5]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3004), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(30)  (.Q (p_nbus_Mem_Alu_R[6]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3005), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(29)  (.Q (p_nbus_Mem_Alu_R[7]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3006), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(28)  (.Q (p_nbus_Mem_Alu_R[8]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3007), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(27)  (.Q (p_nbus_Mem_Alu_R[9]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3008), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(26)  (.Q (p_nbus_Mem_Alu_R[10]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3009), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(25)  (.Q (p_nbus_Mem_Alu_R[11]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3010), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(24)  (.Q (p_nbus_Mem_Alu_R[12]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3011), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(23)  (.Q (p_nbus_Mem_Alu_R[13]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3012), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(22)  (.Q (p_nbus_Mem_Alu_R[14]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3013), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(21)  (.Q (p_nbus_Mem_Alu_R[15]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3014), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(20)  (.Q (p_nbus_Mem_Alu_R[16]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3015), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(19)  (.Q (p_nbus_Mem_Alu_R[17]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3016), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(18)  (.Q (p_nbus_Mem_Alu_R[18]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3017), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(17)  (.Q (p_nbus_Mem_Alu_R[19]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3018), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(16)  (.Q (p_nbus_Mem_Alu_R[20]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3019), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(15)  (.Q (p_nbus_Mem_Alu_R[21]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3020), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(14)  (.Q (p_nbus_Mem_Alu_R[22]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3021), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(13)  (.Q (p_nbus_Mem_Alu_R[23]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3022), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(12)  (.Q (p_nbus_Mem_Alu_R[24]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3023), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(11)  (.Q (p_nbus_Mem_Alu_R[25]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3024), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(10)  (.Q (p_nbus_Mem_Alu_R[26]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3025), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(9)  (.Q (p_nbus_Mem_Alu_R[27]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3026), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(8)  (.Q (p_nbus_Mem_Alu_R[28]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3027), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(7)  (.Q (p_nbus_Mem_Alu_R[29]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3028), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(1)  (.Q (p_nbus_Mem_Alu_R[30]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3029), .R (px3433)) ;
    FDRE \reg_Mem_Alu_R(0)  (.Q (p_nbus_Mem_Alu_R[31]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3030), .R (px3433)) ;
    FDRE \reg_Mem_Rd(2)  (.Q (p_nbus_Mem_Rd[0]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_Rd[0]), .R (px3433)) ;
    FDRE \reg_Mem_Rd(1)  (.Q (p_nbus_Mem_Rd[1]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_Rd[1]), .R (px3433)) ;
    FDRE \reg_Mem_Rd(0)  (.Q (p_nbus_Mem_Rd[2]), .C (p_CLK_int), .CE (p_EN_int)
         , .D (p_nbus_Ex_Rd[2]), .R (px3433)) ;
    FDRE reg_Mem_Wmem (.Q (p_Mem_Wmem), .C (p_CLK_int), .CE (p_EN_int), .D (
         p_Ex_Wmem), .R (px3433)) ;
    FDRE reg_Mem_Reg2reg (.Q (p_Mem_Reg2reg), .C (p_CLK_int), .CE (p_EN_int), .D (
         p_Ex_Reg2reg), .R (px3433)) ;
    FDRE reg_Mem_Wreg (.Q (p_Mem_Wreg), .C (p_CLK_int), .CE (p_EN_int), .D (
         p_Ex_Wreg), .R (px3433)) ;
    LUT6 ix54906z1314 (.O (px3209), .I0 (px3327), .I1 (px3326), .I2 (px3315), .I3 (
         px3314), .I4 (px3309), .I5 (px3308)) ;
         defparam ix54906z1314.INIT = 64'h0000066006600000;
    LUT6 ix55894z1314 (.O (px3210), .I0 (px3336), .I1 (px3335), .I2 (px3321), .I3 (
         px3320), .I4 (px3318), .I5 (px3317)) ;
         defparam ix55894z1314.INIT = 64'h0000066006600000;
    LUT6 ix55895z1314 (.O (px3211), .I0 (px3339), .I1 (px3338), .I2 (px3324), .I3 (
         px3323), .I4 (px3306), .I5 (px3305)) ;
         defparam ix55895z1314.INIT = 64'h0000066006600000;
    LUT6 ix55896z1314 (.O (px3212), .I0 (px3357), .I1 (px3356), .I2 (px3354), .I3 (
         px3353), .I4 (px3330), .I5 (px3329)) ;
         defparam ix55896z1314.INIT = 64'h0000066006600000;
    LUT6 ix55897z1314 (.O (px3213), .I0 (px3363), .I1 (px3362), .I2 (px3360), .I3 (
         px3359), .I4 (px3303), .I5 (px3302)) ;
         defparam ix55897z1314.INIT = 64'h0000066006600000;
    LUT6 ix55898z1314 (.O (px3214), .I0 (px3300), .I1 (px3299), .I2 (px3297), .I3 (
         px3296), .I4 (px3294), .I5 (px3293)) ;
         defparam ix55898z1314.INIT = 64'h0000066006600000;
    LUT6 ix55899z1314 (.O (px3215), .I0 (px3333), .I1 (px3332), .I2 (px3291), .I3 (
         px3290), .I4 (px3288), .I5 (px3287)) ;
         defparam ix55899z1314.INIT = 64'h0000066006600000;
    LUT6 ix59885z1318 (.O (px3253), .I0 (px3255), .I1 (nx59885z3), .I2 (
         \p_Rs_1_0(2)  ), .I3 (\p_Rs_1_0(0)  ), .I4 (p_nbus_Mem_Rd[0]), .I5 (
         p_nbus_Mem_Rd[2])) ;
         defparam ix59885z1318.INIT = 64'h4000040000400004;
    LUT5 ix59885z1315 (.O (nx59885z3), .I0 (\p_Rs_1_0(1)  ), .I1 (
         p_nbus_Mem_Rd[0]), .I2 (p_nbus_Mem_Rd[1]), .I3 (p_nbus_Mem_Rd[2]), .I4 (
         p_Mem_Wreg)) ;
         defparam ix59885z1315.INIT = 32'hA5A40000;
    LUT6 ix59888z1314 (.O (px3256), .I0 (px3258), .I1 (nx59888z3), .I2 (
         p_nbus_Mem_Rd[0]), .I3 (p_nbus_Mem_Rd[1]), .I4 (p_nbus_Mem_Rd[2]), .I5 (
         p_Mem_Wreg)) ;
         defparam ix59888z1314.INIT = 64'h4444444000000000;
    LUT6 ix59888z1828 (.O (nx59888z3), .I0 (\p_Rt_1_0(2)  ), .I1 (\p_Rt_1_0(1)  
         ), .I2 (\p_Rt_1_0(0)  ), .I3 (p_nbus_Mem_Rd[0]), .I4 (p_nbus_Mem_Rd[1])
         , .I5 (p_nbus_Mem_Rd[2])) ;
         defparam ix59888z1828.INIT = 64'h8040201008040201;
    LUT5 ix62880z5205 (.O (px3287), .I0 (px3487), .I1 (p_nbus_Ex_D1[5]), .I2 (
         p_nbus_Mem_Alu_R[5]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix62880z5205.INIT = 32'h33AA0F33;
    LUT5 ix63870z5205 (.O (px3290), .I0 (px3486), .I1 (p_nbus_Ex_D1[6]), .I2 (
         p_nbus_Mem_Alu_R[6]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix63870z5205.INIT = 32'h33AA0F33;
    LUT5 ix63873z5205 (.O (px3293), .I0 (px3485), .I1 (p_nbus_Ex_D1[7]), .I2 (
         p_nbus_Mem_Alu_R[7]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix63873z5205.INIT = 32'h33AA0F33;
    LUT5 ix63876z5205 (.O (px3296), .I0 (px3484), .I1 (p_nbus_Ex_D1[8]), .I2 (
         p_nbus_Mem_Alu_R[8]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix63876z5205.INIT = 32'h33AA0F33;
    LUT5 ix63879z5205 (.O (px3299), .I0 (px3483), .I1 (p_nbus_Ex_D1[9]), .I2 (
         p_nbus_Mem_Alu_R[9]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix63879z5205.INIT = 32'h33AA0F33;
    LUT5 ix332z5205 (.O (px3302), .I0 (px3482), .I1 (p_nbus_Ex_D1[10]), .I2 (
         p_nbus_Mem_Alu_R[10]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix332z5205.INIT = 32'h33AA0F33;
    LUT5 ix335z5205 (.O (px3305), .I0 (px3481), .I1 (p_nbus_Ex_D1[11]), .I2 (
         p_nbus_Mem_Alu_R[11]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix335z5205.INIT = 32'h33AA0F33;
    LUT5 ix338z5205 (.O (px3308), .I0 (px3480), .I1 (p_nbus_Ex_D1[12]), .I2 (
         p_nbus_Mem_Alu_R[12]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix338z5205.INIT = 32'h33AA0F33;
    LUT5 ix1328z5205 (.O (px3311), .I0 (px3479), .I1 (p_nbus_Ex_D1[13]), .I2 (
         p_nbus_Mem_Alu_R[13]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix1328z5205.INIT = 32'h33AA0F33;
    LUT5 ix1331z5205 (.O (px3314), .I0 (px3478), .I1 (p_nbus_Ex_D1[14]), .I2 (
         p_nbus_Mem_Alu_R[14]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix1331z5205.INIT = 32'h33AA0F33;
    LUT5 ix1334z5205 (.O (px3317), .I0 (px3477), .I1 (p_nbus_Ex_D1[15]), .I2 (
         p_nbus_Mem_Alu_R[15]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix1334z5205.INIT = 32'h33AA0F33;
    LUT5 ix2324z5205 (.O (px3320), .I0 (px3476), .I1 (p_nbus_Ex_D1[16]), .I2 (
         p_nbus_Mem_Alu_R[16]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix2324z5205.INIT = 32'h33AA0F33;
    LUT5 ix2327z5205 (.O (px3323), .I0 (px3475), .I1 (p_nbus_Ex_D1[17]), .I2 (
         p_nbus_Mem_Alu_R[17]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix2327z5205.INIT = 32'h33AA0F33;
    LUT5 ix2330z5205 (.O (px3326), .I0 (px3474), .I1 (p_nbus_Ex_D1[18]), .I2 (
         p_nbus_Mem_Alu_R[18]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix2330z5205.INIT = 32'h33AA0F33;
    LUT5 ix2333z5205 (.O (px3329), .I0 (px3473), .I1 (p_nbus_Ex_D1[19]), .I2 (
         p_nbus_Mem_Alu_R[19]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix2333z5205.INIT = 32'h33AA0F33;
    LUT5 ix3323z5205 (.O (px3332), .I0 (px3472), .I1 (p_nbus_Ex_D1[20]), .I2 (
         p_nbus_Mem_Alu_R[20]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix3323z5205.INIT = 32'h33AA0F33;
    LUT5 ix3326z5205 (.O (px3335), .I0 (px3471), .I1 (p_nbus_Ex_D1[21]), .I2 (
         p_nbus_Mem_Alu_R[21]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix3326z5205.INIT = 32'h33AA0F33;
    LUT5 ix3329z5205 (.O (px3338), .I0 (px3470), .I1 (p_nbus_Ex_D1[22]), .I2 (
         p_nbus_Mem_Alu_R[22]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix3329z5205.INIT = 32'h33AA0F33;
    LUT5 ix4319z5205 (.O (px3341), .I0 (px3469), .I1 (p_nbus_Ex_D1[23]), .I2 (
         p_nbus_Mem_Alu_R[23]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix4319z5205.INIT = 32'h33AA0F33;
    LUT5 ix4323z5205 (.O (px3345), .I0 (px3468), .I1 (p_nbus_Ex_D1[24]), .I2 (
         p_nbus_Mem_Alu_R[24]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix4323z5205.INIT = 32'h33AA0F33;
    LUT6 ix4325z1313 (.O (px3347), .I0 (p_nbus_Mem_Alu_R[24]), .I1 (
         p_nbus_Wb_D[29]), .I2 (p_nbus_Wb_Alu_R[29]), .I3 (p_Wb_Reg2reg), .I4 (
         p_nbus_Ex_Fwd_B[0]), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix4325z1313.INIT = 64'hFFFF0F335555FFFF;
    LUT5 ix4327z5205 (.O (px3349), .I0 (px3467), .I1 (p_nbus_Ex_D1[25]), .I2 (
         p_nbus_Mem_Alu_R[25]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix4327z5205.INIT = 32'h33AA0F33;
    LUT6 ix5316z1313 (.O (px3351), .I0 (p_nbus_Mem_Alu_R[25]), .I1 (
         p_nbus_Wb_D[30]), .I2 (p_nbus_Wb_Alu_R[30]), .I3 (p_Wb_Reg2reg), .I4 (
         p_nbus_Ex_Fwd_B[0]), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix5316z1313.INIT = 64'hFFFF0F335555FFFF;
    LUT5 ix5318z5205 (.O (px3353), .I0 (px3466), .I1 (p_nbus_Ex_D1[26]), .I2 (
         p_nbus_Mem_Alu_R[26]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix5318z5205.INIT = 32'h33AA0F33;
    LUT5 ix5321z5205 (.O (px3356), .I0 (px3465), .I1 (p_nbus_Ex_D1[27]), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix5321z5205.INIT = 32'h33AA0F33;
    LUT5 ix5324z5205 (.O (px3359), .I0 (px3464), .I1 (p_nbus_Ex_D1[28]), .I2 (
         p_nbus_Mem_Alu_R[28]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix5324z5205.INIT = 32'h33AA0F33;
    LUT5 ix6314z5205 (.O (px3362), .I0 (px3463), .I1 (p_nbus_Ex_D1[29]), .I2 (
         p_nbus_Mem_Alu_R[29]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix6314z5205.INIT = 32'h33AA0F33;
    LUT5 ix6317z5205 (.O (px3365), .I0 (px3457), .I1 (p_nbus_Ex_D1[30]), .I2 (
         p_nbus_Mem_Alu_R[30]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix6317z5205.INIT = 32'h33AA0F33;
    LUT6 ix6319z1313 (.O (px3367), .I0 (p_nbus_Mem_Alu_R[30]), .I1 (
         p_nbus_Wb_D[31]), .I2 (p_nbus_Wb_Alu_R[31]), .I3 (p_Wb_Reg2reg), .I4 (
         p_nbus_Ex_Fwd_B[0]), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix6319z1313.INIT = 64'hFFFF0F335555FFFF;
    LUT6 ix6320z25687 (.O (px3368), .I0 (p_nbus_Ex_D1[31]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (p_nbus_Ex_Aluc[0]), .I5 (px3373)) ;
         defparam ix6320z25687.INIT = 64'h0000000000005F35;
    LUT2 ix24571z1316 (.O (px3433), .I0 (p_EN_int), .I1 (p_CLR_N_int)) ;
         defparam ix24571z1316.INIT = 4'h2;
    LUT3 ix14295z1334 (.O (px3435), .I0 (p_nbus_Ex_Aluc[1]), .I1 (
         p_nbus_Ex_Aluc[2]), .I2 (p_nbus_Ex_Aluc[0])) ;
         defparam ix14295z1334.INIT = 8'h14;
    LUT2 ix14296z1318 (.O (px3436), .I0 (p_nbus_Ex_Aluc[1]), .I1 (
         p_nbus_Ex_Aluc[0])) ;
         defparam ix14296z1318.INIT = 4'h4;
endmodule


module ALU_0 ( p_nbus_Wb_Alu_R, p_nbus_Wb_D, p_nbus_Ex_D2, \p_Ex_Op(0)  , px3439, 
               px3432, px3428, px3424, px3420, p_nbus_Ex_D1, p_nbus_Ex_Aluc, 
               p_nbus_Mem_Alu_R, \p_Ex_Extimm(13)  , px3343, p_nbus_Ex_Fwd_B, 
               px3041, px3430, px3040, px3426, px3039, px3422, px3038, px3037, 
               px3368, px3369, px3030, px3365, px3029, px3362, px3028, px3359, 
               px3027, px3356, px3026, px3353, px3025, px3349, px3024, px3345, 
               px3023, px3341, px3022, px3338, px3021, px3335, px3020, px3332, 
               px3019, px3329, px3018, px3326, px3017, px3323, px3016, px3320, 
               px3015, px3317, px3014, px3314, px3013, px3311, px3012, px3308, 
               px3011, px3305, px3010, px3302, px3009, px3299, px3008, px3296, 
               px3007, px3293, px3006, px3290, px3005, px3435, px3436, px3287, 
               px3004, p_Wb_Reg2reg, p_Ex_Aluqb, \p_Ex_Extimm(0)  , px3370, 
               px3371, px3373, px3366, px3457, px3419, px3423, px3427, px3431, 
               px3462, px3363, px3463, px3360, px3464, px3357, px3465, px3354, 
               px3466, px3350, px3467, px3346, px3468, px3469, px3339, px3470, 
               px3336, px3471, px3333, px3472, px3330, px3473, px3327, px3474, 
               px3324, px3475, px3321, px3476, px3318, px3477, px3315, px3478, 
               px3312, px3479, px3309, px3480, px3306, px3481, px3303, px3482, 
               px3300, px3483, px3297, px3484, px3294, px3485, px3291, px3486, 
               px3288, px3487, p_nbus_Ex_Fwd_A, px2963, p_Ex_Z, px3206, px3209, 
               px3210, px3211, px3212, px3213, px3214, px3215, px2855, px2964, 
               px2965, px2966, px2967, px2968, px2969, px2970, px2971, px2972, 
               px2973, px2974, px2975, px2976, px2977, px2978, px2979, px2980, 
               px2981, px2982, px2983, px2984, px2985, px2986, px2987, px2988, 
               px2989, px2990, px2991, px2992, px2993, px2994, px2857 ) ;

    input [31:0]p_nbus_Wb_Alu_R ;
    input [31:0]p_nbus_Wb_D ;
    input [31:6]p_nbus_Ex_D2 ;
    input \p_Ex_Op(0)   ;
    output px3439 ;
    output px3432 ;
    output px3428 ;
    output px3424 ;
    output px3420 ;
    input [31:0]p_nbus_Ex_D1 ;
    input [2:0]p_nbus_Ex_Aluc ;
    input [31:0]p_nbus_Mem_Alu_R ;
    input \p_Ex_Extimm(13)   ;
    output px3343 ;
    input [1:0]p_nbus_Ex_Fwd_B ;
    output px3041 ;
    output px3430 ;
    output px3040 ;
    output px3426 ;
    output px3039 ;
    output px3422 ;
    output px3038 ;
    output px3037 ;
    input px3368 ;
    input px3369 ;
    output px3030 ;
    input px3365 ;
    output px3029 ;
    input px3362 ;
    output px3028 ;
    input px3359 ;
    output px3027 ;
    input px3356 ;
    output px3026 ;
    input px3353 ;
    output px3025 ;
    input px3349 ;
    output px3024 ;
    input px3345 ;
    output px3023 ;
    input px3341 ;
    output px3022 ;
    input px3338 ;
    output px3021 ;
    input px3335 ;
    output px3020 ;
    input px3332 ;
    output px3019 ;
    input px3329 ;
    output px3018 ;
    input px3326 ;
    output px3017 ;
    input px3323 ;
    output px3016 ;
    input px3320 ;
    output px3015 ;
    input px3317 ;
    output px3014 ;
    input px3314 ;
    output px3013 ;
    input px3311 ;
    output px3012 ;
    input px3308 ;
    output px3011 ;
    input px3305 ;
    output px3010 ;
    input px3302 ;
    output px3009 ;
    input px3299 ;
    output px3008 ;
    input px3296 ;
    output px3007 ;
    input px3293 ;
    output px3006 ;
    input px3290 ;
    output px3005 ;
    input px3435 ;
    input px3436 ;
    input px3287 ;
    output px3004 ;
    input p_Wb_Reg2reg ;
    input p_Ex_Aluqb ;
    input \p_Ex_Extimm(0)   ;
    output px3370 ;
    output px3371 ;
    output px3373 ;
    input px3366 ;
    output px3457 ;
    input px3419 ;
    input px3423 ;
    input px3427 ;
    output px3431 ;
    output px3462 ;
    output px3363 ;
    output px3463 ;
    output px3360 ;
    output px3464 ;
    output px3357 ;
    output px3465 ;
    output px3354 ;
    output px3466 ;
    input px3350 ;
    output px3467 ;
    input px3346 ;
    output px3468 ;
    output px3469 ;
    output px3339 ;
    output px3470 ;
    output px3336 ;
    output px3471 ;
    output px3333 ;
    output px3472 ;
    output px3330 ;
    output px3473 ;
    output px3327 ;
    output px3474 ;
    output px3324 ;
    output px3475 ;
    output px3321 ;
    output px3476 ;
    output px3318 ;
    output px3477 ;
    output px3315 ;
    output px3478 ;
    output px3312 ;
    output px3479 ;
    output px3309 ;
    output px3480 ;
    output px3306 ;
    output px3481 ;
    output px3303 ;
    output px3482 ;
    output px3300 ;
    output px3483 ;
    output px3297 ;
    output px3484 ;
    output px3294 ;
    output px3485 ;
    output px3291 ;
    output px3486 ;
    output px3288 ;
    output px3487 ;
    input [1:0]p_nbus_Ex_Fwd_A ;
    output px2963 ;
    output p_Ex_Z ;
    input px3206 ;
    input px3209 ;
    input px3210 ;
    input px3211 ;
    input px3212 ;
    input px3213 ;
    input px3214 ;
    input px3215 ;
    input px2855 ;
    output px2964 ;
    output px2965 ;
    output px2966 ;
    output px2967 ;
    output px2968 ;
    output px2969 ;
    output px2970 ;
    output px2971 ;
    output px2972 ;
    output px2973 ;
    output px2974 ;
    output px2975 ;
    output px2976 ;
    output px2977 ;
    output px2978 ;
    output px2979 ;
    output px2980 ;
    output px2981 ;
    output px2982 ;
    output px2983 ;
    output px2984 ;
    output px2985 ;
    output px2986 ;
    output px2987 ;
    output px2988 ;
    output px2989 ;
    output px2990 ;
    output px2991 ;
    output px2992 ;
    output px2993 ;
    output px2994 ;
    input px2857 ;

    wire nx36948z7, nx36948z4, nx36947z2, nx35959z2, nx35958z2, nx35957z3, 
         nx35957z2, nx35950z2, nx34962z3, nx34961z3, nx34960z3, nx34959z3, 
         nx34958z3, nx34957z3, nx34956z3, nx34955z3, nx34954z3, nx34953z3, 
         nx33965z3, nx33964z3, nx33963z3, nx33962z3, nx33961z3, nx33960z3, 
         nx33959z3, nx33958z3, nx33957z3, nx33956z3, nx32968z3, nx32967z3, 
         nx32966z3, nx32965z3, nx32964z3, nx32963z3, nx20404z3, nx20406z3, 
         nx20407z3, nx20408z3, nx20409z3, nx36948z2, nx321z5, nx35950z5, 
         nx2313z4;
    wire [31:0]alu_R_0n0s6;
    wire nx2313z1, nx2312z4, nx2312z1, nx1324z4, nx1324z1, nx1323z4, nx1323z1, 
         nx1322z4, nx1322z1, nx1321z4, nx1321z1, nx1320z4, nx1320z1, nx1319z4, 
         nx1319z1, nx1318z4, nx1318z1, nx1317z4, nx1317z1, nx1316z4, nx1316z1, 
         nx1315z4, nx1315z1, nx327z4, nx327z1, nx326z4, nx326z1, nx325z4, 
         nx325z1, nx324z4, nx324z1, nx323z4, nx323z1, nx322z4, nx322z1, nx321z4, 
         nx321z1, nx320z4, nx320z1, nx319z4, nx319z1, nx318z4, nx318z1, 
         nx63490z4, nx63490z1, nx63491z4, nx63491z1, nx63492z4, nx63492z1, 
         nx58118z2, nx58118z1, nx63494z2, nx63494z1, nx63495z2, nx63495z1, 
         nx63496z2, nx63496z1, nx63497z2, nx63497z1, nx63498z2, nx63498z1, 
         nx63499z2, nx60029z21, nx60029z1, nx60029z19, nx60029z2, nx60029z18, 
         nx60029z3, nx60029z4, nx60029z5, nx60029z6, nx60029z7, nx60029z8, 
         nx60029z9, nx60029z10, nx14591z2;
    wire [31:0]alu_R_0n0s3;
    wire nx14591z1, nx14590z2, nx14590z1, nx13602z2, nx13602z1, nx13601z2, 
         nx13601z1, nx13600z2, nx13600z1, nx13599z2, nx13599z1, nx13598z2, 
         nx13598z1, nx13597z2, nx13597z1, nx13596z2, nx13596z1, nx13595z2, 
         nx13595z1, nx13594z2, nx13594z1, nx13593z2, nx13593z1, nx12605z2, 
         nx12605z1, nx12604z2, nx12604z1, nx12603z2, nx12603z1, nx12602z2, 
         nx12602z1, nx12601z2, nx12601z1, nx12600z2, nx12600z1, nx12599z2, 
         nx12599z1, nx12598z2, nx12598z1, nx12597z2, nx12597z1, nx12596z2, 
         nx12596z1, nx39748z2, nx39748z1, nx39749z2, nx39749z1, nx39750z2, 
         nx39750z1, nx39751z2, nx39751z1, nx20409z4, nx20409z1, nx20408z4, 
         nx20408z1, nx20407z4, nx20407z1, nx20406z4, nx20406z1, nx20405z4, 
         nx20405z1, nx20404z4;



    XORCY R_add32_0i1_xorcy_0 (.O (alu_R_0n0s3[0]), .CI (px2857), .LI (nx20404z4
          )) ;
    XORCY R_add32_0i1_xorcy_1 (.O (alu_R_0n0s3[1]), .CI (nx20405z1), .LI (
          nx20405z4)) ;
    XORCY R_add32_0i1_xorcy_2 (.O (alu_R_0n0s3[2]), .CI (nx20406z1), .LI (
          nx20406z4)) ;
    XORCY R_add32_0i1_xorcy_3 (.O (alu_R_0n0s3[3]), .CI (nx20407z1), .LI (
          nx20407z4)) ;
    XORCY R_add32_0i1_xorcy_4 (.O (alu_R_0n0s3[4]), .CI (nx20408z1), .LI (
          nx20408z4)) ;
    XORCY R_add32_0i1_xorcy_5 (.O (alu_R_0n0s3[5]), .CI (nx20409z1), .LI (
          nx20409z4)) ;
    XORCY R_add32_0i1_xorcy_6 (.O (alu_R_0n0s3[6]), .CI (nx39751z1), .LI (
          nx39751z2)) ;
    XORCY R_add32_0i1_xorcy_7 (.O (alu_R_0n0s3[7]), .CI (nx39750z1), .LI (
          nx39750z2)) ;
    XORCY R_add32_0i1_xorcy_8 (.O (alu_R_0n0s3[8]), .CI (nx39749z1), .LI (
          nx39749z2)) ;
    XORCY R_add32_0i1_xorcy_9 (.O (alu_R_0n0s3[9]), .CI (nx39748z1), .LI (
          nx39748z2)) ;
    XORCY R_add32_0i1_xorcy_10 (.O (alu_R_0n0s3[10]), .CI (nx12596z1), .LI (
          nx12596z2)) ;
    XORCY R_add32_0i1_xorcy_11 (.O (alu_R_0n0s3[11]), .CI (nx12597z1), .LI (
          nx12597z2)) ;
    XORCY R_add32_0i1_xorcy_12 (.O (alu_R_0n0s3[12]), .CI (nx12598z1), .LI (
          nx12598z2)) ;
    XORCY R_add32_0i1_xorcy_13 (.O (alu_R_0n0s3[13]), .CI (nx12599z1), .LI (
          nx12599z2)) ;
    XORCY R_add32_0i1_xorcy_14 (.O (alu_R_0n0s3[14]), .CI (nx12600z1), .LI (
          nx12600z2)) ;
    XORCY R_add32_0i1_xorcy_15 (.O (alu_R_0n0s3[15]), .CI (nx12601z1), .LI (
          nx12601z2)) ;
    XORCY R_add32_0i1_xorcy_16 (.O (alu_R_0n0s3[16]), .CI (nx12602z1), .LI (
          nx12602z2)) ;
    XORCY R_add32_0i1_xorcy_17 (.O (alu_R_0n0s3[17]), .CI (nx12603z1), .LI (
          nx12603z2)) ;
    XORCY R_add32_0i1_xorcy_18 (.O (alu_R_0n0s3[18]), .CI (nx12604z1), .LI (
          nx12604z2)) ;
    XORCY R_add32_0i1_xorcy_19 (.O (alu_R_0n0s3[19]), .CI (nx12605z1), .LI (
          nx12605z2)) ;
    XORCY R_add32_0i1_xorcy_20 (.O (alu_R_0n0s3[20]), .CI (nx13593z1), .LI (
          nx13593z2)) ;
    XORCY R_add32_0i1_xorcy_21 (.O (alu_R_0n0s3[21]), .CI (nx13594z1), .LI (
          nx13594z2)) ;
    XORCY R_add32_0i1_xorcy_22 (.O (alu_R_0n0s3[22]), .CI (nx13595z1), .LI (
          nx13595z2)) ;
    XORCY R_add32_0i1_xorcy_23 (.O (alu_R_0n0s3[23]), .CI (nx13596z1), .LI (
          nx13596z2)) ;
    XORCY R_add32_0i1_xorcy_24 (.O (alu_R_0n0s3[24]), .CI (nx13597z1), .LI (
          nx13597z2)) ;
    XORCY R_add32_0i1_xorcy_25 (.O (alu_R_0n0s3[25]), .CI (nx13598z1), .LI (
          nx13598z2)) ;
    XORCY R_add32_0i1_xorcy_26 (.O (alu_R_0n0s3[26]), .CI (nx13599z1), .LI (
          nx13599z2)) ;
    XORCY R_add32_0i1_xorcy_27 (.O (alu_R_0n0s3[27]), .CI (nx13600z1), .LI (
          nx13600z2)) ;
    XORCY R_add32_0i1_xorcy_28 (.O (alu_R_0n0s3[28]), .CI (nx13601z1), .LI (
          nx13601z2)) ;
    XORCY R_add32_0i1_xorcy_29 (.O (alu_R_0n0s3[29]), .CI (nx13602z1), .LI (
          nx13602z2)) ;
    XORCY R_add32_0i1_xorcy_30 (.O (alu_R_0n0s3[30]), .CI (nx14590z1), .LI (
          nx14590z2)) ;
    XORCY R_add32_0i1_xorcy_31 (.O (alu_R_0n0s3[31]), .CI (nx14591z1), .LI (
          nx14591z2)) ;
    MUXCY Z_eq_0_ix60029z52223 (.O (p_Ex_Z), .CI (nx60029z1), .DI (px2857), .S (
          nx60029z21)) ;
    XORCY R_sub32_0i5_xorcy_0 (.O (alu_R_0n0s6[0]), .CI (px2855), .LI (nx63499z2
          )) ;
    XORCY R_sub32_0i5_xorcy_1 (.O (alu_R_0n0s6[1]), .CI (nx63498z1), .LI (
          nx63498z2)) ;
    XORCY R_sub32_0i5_xorcy_2 (.O (alu_R_0n0s6[2]), .CI (nx63497z1), .LI (
          nx63497z2)) ;
    XORCY R_sub32_0i5_xorcy_3 (.O (alu_R_0n0s6[3]), .CI (nx63496z1), .LI (
          nx63496z2)) ;
    XORCY R_sub32_0i5_xorcy_4 (.O (alu_R_0n0s6[4]), .CI (nx63495z1), .LI (
          nx63495z2)) ;
    XORCY R_sub32_0i5_xorcy_5 (.O (alu_R_0n0s6[5]), .CI (nx63494z1), .LI (
          nx63494z2)) ;
    XORCY R_sub32_0i5_xorcy_6 (.O (alu_R_0n0s6[6]), .CI (nx58118z1), .LI (
          nx58118z2)) ;
    XORCY R_sub32_0i5_xorcy_7 (.O (alu_R_0n0s6[7]), .CI (nx63492z1), .LI (
          nx63492z4)) ;
    XORCY R_sub32_0i5_xorcy_8 (.O (alu_R_0n0s6[8]), .CI (nx63491z1), .LI (
          nx63491z4)) ;
    XORCY R_sub32_0i5_xorcy_9 (.O (alu_R_0n0s6[9]), .CI (nx63490z1), .LI (
          nx63490z4)) ;
    XORCY R_sub32_0i5_xorcy_10 (.O (alu_R_0n0s6[10]), .CI (nx318z1), .LI (
          nx318z4)) ;
    XORCY R_sub32_0i5_xorcy_11 (.O (alu_R_0n0s6[11]), .CI (nx319z1), .LI (
          nx319z4)) ;
    XORCY R_sub32_0i5_xorcy_12 (.O (alu_R_0n0s6[12]), .CI (nx320z1), .LI (
          nx320z4)) ;
    XORCY R_sub32_0i5_xorcy_13 (.O (alu_R_0n0s6[13]), .CI (nx321z1), .LI (
          nx321z4)) ;
    XORCY R_sub32_0i5_xorcy_14 (.O (alu_R_0n0s6[14]), .CI (nx322z1), .LI (
          nx322z4)) ;
    XORCY R_sub32_0i5_xorcy_15 (.O (alu_R_0n0s6[15]), .CI (nx323z1), .LI (
          nx323z4)) ;
    XORCY R_sub32_0i5_xorcy_16 (.O (alu_R_0n0s6[16]), .CI (nx324z1), .LI (
          nx324z4)) ;
    XORCY R_sub32_0i5_xorcy_17 (.O (alu_R_0n0s6[17]), .CI (nx325z1), .LI (
          nx325z4)) ;
    XORCY R_sub32_0i5_xorcy_18 (.O (alu_R_0n0s6[18]), .CI (nx326z1), .LI (
          nx326z4)) ;
    XORCY R_sub32_0i5_xorcy_19 (.O (alu_R_0n0s6[19]), .CI (nx327z1), .LI (
          nx327z4)) ;
    XORCY R_sub32_0i5_xorcy_20 (.O (alu_R_0n0s6[20]), .CI (nx1315z1), .LI (
          nx1315z4)) ;
    XORCY R_sub32_0i5_xorcy_21 (.O (alu_R_0n0s6[21]), .CI (nx1316z1), .LI (
          nx1316z4)) ;
    XORCY R_sub32_0i5_xorcy_22 (.O (alu_R_0n0s6[22]), .CI (nx1317z1), .LI (
          nx1317z4)) ;
    XORCY R_sub32_0i5_xorcy_23 (.O (alu_R_0n0s6[23]), .CI (nx1318z1), .LI (
          nx1318z4)) ;
    XORCY R_sub32_0i5_xorcy_24 (.O (alu_R_0n0s6[24]), .CI (nx1319z1), .LI (
          nx1319z4)) ;
    XORCY R_sub32_0i5_xorcy_25 (.O (alu_R_0n0s6[25]), .CI (nx1320z1), .LI (
          nx1320z4)) ;
    XORCY R_sub32_0i5_xorcy_26 (.O (alu_R_0n0s6[26]), .CI (nx1321z1), .LI (
          nx1321z4)) ;
    XORCY R_sub32_0i5_xorcy_27 (.O (alu_R_0n0s6[27]), .CI (nx1322z1), .LI (
          nx1322z4)) ;
    XORCY R_sub32_0i5_xorcy_28 (.O (alu_R_0n0s6[28]), .CI (nx1323z1), .LI (
          nx1323z4)) ;
    XORCY R_sub32_0i5_xorcy_29 (.O (alu_R_0n0s6[29]), .CI (nx1324z1), .LI (
          nx1324z4)) ;
    XORCY R_sub32_0i5_xorcy_30 (.O (alu_R_0n0s6[30]), .CI (nx2312z1), .LI (
          nx2312z4)) ;
    XORCY R_sub32_0i5_xorcy_31 (.O (alu_R_0n0s6[31]), .CI (nx2313z1), .LI (
          nx2313z4)) ;
    MUXCY R_sub32_0i5_muxcy_31 (.O (nx35950z5), .CI (nx2313z1), .DI (px2963), .S (
          nx2313z4)) ;
    LUT6 ix2313z21849 (.O (nx2313z4), .I0 (p_nbus_Ex_D1[0]), .I1 (
         p_nbus_Mem_Alu_R[0]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3487), .I5 (px3288)) ;
         defparam ix2313z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix2312z21849 (.O (nx2312z4), .I0 (p_nbus_Ex_D1[1]), .I1 (
         p_nbus_Mem_Alu_R[1]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3486), .I5 (px3291)) ;
         defparam ix2312z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1324z21849 (.O (nx1324z4), .I0 (p_nbus_Ex_D1[2]), .I1 (
         p_nbus_Mem_Alu_R[2]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3485), .I5 (px3294)) ;
         defparam ix1324z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1323z21849 (.O (nx1323z4), .I0 (p_nbus_Ex_D1[3]), .I1 (
         p_nbus_Mem_Alu_R[3]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3484), .I5 (px3297)) ;
         defparam ix1323z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1322z21849 (.O (nx1322z4), .I0 (p_nbus_Ex_D1[4]), .I1 (
         p_nbus_Mem_Alu_R[4]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3483), .I5 (px3300)) ;
         defparam ix1322z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1321z21849 (.O (nx1321z4), .I0 (p_nbus_Ex_D1[5]), .I1 (
         p_nbus_Mem_Alu_R[5]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3482), .I5 (px3303)) ;
         defparam ix1321z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1320z21849 (.O (nx1320z4), .I0 (p_nbus_Ex_D1[6]), .I1 (
         p_nbus_Mem_Alu_R[6]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3481), .I5 (px3306)) ;
         defparam ix1320z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1319z21849 (.O (nx1319z4), .I0 (p_nbus_Ex_D1[7]), .I1 (
         p_nbus_Mem_Alu_R[7]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3480), .I5 (px3309)) ;
         defparam ix1319z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1318z21849 (.O (nx1318z4), .I0 (p_nbus_Ex_D1[8]), .I1 (
         p_nbus_Mem_Alu_R[8]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3479), .I5 (px3312)) ;
         defparam ix1318z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1317z21849 (.O (nx1317z4), .I0 (p_nbus_Ex_D1[9]), .I1 (
         p_nbus_Mem_Alu_R[9]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3478), .I5 (px3315)) ;
         defparam ix1317z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1316z21849 (.O (nx1316z4), .I0 (p_nbus_Ex_D1[10]), .I1 (
         p_nbus_Mem_Alu_R[10]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3477), .I5 (px3318)) ;
         defparam ix1316z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix1315z21849 (.O (nx1315z4), .I0 (p_nbus_Ex_D1[11]), .I1 (
         p_nbus_Mem_Alu_R[11]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3476), .I5 (px3321)) ;
         defparam ix1315z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix327z21849 (.O (nx327z4), .I0 (p_nbus_Ex_D1[12]), .I1 (
         p_nbus_Mem_Alu_R[12]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3475), .I5 (px3324)) ;
         defparam ix327z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix326z21849 (.O (nx326z4), .I0 (p_nbus_Ex_D1[13]), .I1 (
         p_nbus_Mem_Alu_R[13]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3474), .I5 (px3327)) ;
         defparam ix326z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix325z21849 (.O (nx325z4), .I0 (p_nbus_Ex_D1[14]), .I1 (
         p_nbus_Mem_Alu_R[14]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3473), .I5 (px3330)) ;
         defparam ix325z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix324z21849 (.O (nx324z4), .I0 (p_nbus_Ex_D1[15]), .I1 (
         p_nbus_Mem_Alu_R[15]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3472), .I5 (px3333)) ;
         defparam ix324z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix323z21849 (.O (nx323z4), .I0 (p_nbus_Ex_D1[16]), .I1 (
         p_nbus_Mem_Alu_R[16]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3471), .I5 (px3336)) ;
         defparam ix323z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix322z21849 (.O (nx322z4), .I0 (p_nbus_Ex_D1[17]), .I1 (
         p_nbus_Mem_Alu_R[17]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3470), .I5 (px3339)) ;
         defparam ix322z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix321z46318 (.O (nx321z4), .I0 (p_nbus_Ex_D1[18]), .I1 (
         p_nbus_Mem_Alu_R[18]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3469), .I5 (nx321z5)) ;
         defparam ix321z46318.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix320z46318 (.O (nx320z4), .I0 (p_nbus_Ex_D1[19]), .I1 (
         p_nbus_Mem_Alu_R[19]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3468), .I5 (px3346)) ;
         defparam ix320z46318.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix319z46318 (.O (nx319z4), .I0 (p_nbus_Ex_D1[20]), .I1 (
         p_nbus_Mem_Alu_R[20]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3467), .I5 (px3350)) ;
         defparam ix319z46318.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix318z21849 (.O (nx318z4), .I0 (p_nbus_Ex_D1[21]), .I1 (
         p_nbus_Mem_Alu_R[21]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3466), .I5 (px3354)) ;
         defparam ix318z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix63490z21849 (.O (nx63490z4), .I0 (p_nbus_Ex_D1[22]), .I1 (
         p_nbus_Mem_Alu_R[22]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3465), .I5 (px3357)) ;
         defparam ix63490z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix63491z21849 (.O (nx63491z4), .I0 (p_nbus_Ex_D1[23]), .I1 (
         p_nbus_Mem_Alu_R[23]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3464), .I5 (px3360)) ;
         defparam ix63491z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix63492z21849 (.O (nx63492z4), .I0 (p_nbus_Ex_D1[24]), .I1 (
         p_nbus_Mem_Alu_R[24]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3463), .I5 (px3363)) ;
         defparam ix63492z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix58118z46316 (.O (nx58118z2), .I0 (p_nbus_Ex_D1[25]), .I1 (
         p_nbus_Mem_Alu_R[25]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3462), .I5 (nx36948z2)) ;
         defparam ix58118z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix63494z46316 (.O (nx63494z2), .I0 (p_nbus_Ex_D1[26]), .I1 (
         p_nbus_Mem_Alu_R[26]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20409z3), .I5 (px3431)) ;
         defparam ix63494z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix63495z46316 (.O (nx63495z2), .I0 (p_nbus_Ex_D1[27]), .I1 (
         p_nbus_Mem_Alu_R[27]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20408z3), .I5 (px3427)) ;
         defparam ix63495z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix63496z46316 (.O (nx63496z2), .I0 (p_nbus_Ex_D1[28]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20407z3), .I5 (px3423)) ;
         defparam ix63496z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix63497z46316 (.O (nx63497z2), .I0 (p_nbus_Ex_D1[29]), .I1 (
         p_nbus_Mem_Alu_R[29]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20406z3), .I5 (px3419)) ;
         defparam ix63497z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix63498z46316 (.O (nx63498z2), .I0 (p_nbus_Ex_D1[30]), .I1 (
         p_nbus_Mem_Alu_R[30]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3457), .I5 (px3366)) ;
         defparam ix63498z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix20404z58113 (.O (nx20404z4), .I0 (nx20404z3), .I1 (px3373), .I2 (
         px3371), .I3 (px3370), .I4 (\p_Ex_Extimm(0)  ), .I5 (p_Ex_Aluqb)) ;
         defparam ix20404z58113.INIT = 64'h22D222D22222DDDD;
    LUT5 ix2313z62958 (.O (px2963), .I0 (px3487), .I1 (p_nbus_Ex_D1[0]), .I2 (
         p_nbus_Mem_Alu_R[0]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix2313z62958.INIT = 32'hCC55F0CC;
    LUT5 ix2312z62958 (.O (px2964), .I0 (px3486), .I1 (p_nbus_Ex_D1[1]), .I2 (
         p_nbus_Mem_Alu_R[1]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix2312z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1324z62958 (.O (px2965), .I0 (px3485), .I1 (p_nbus_Ex_D1[2]), .I2 (
         p_nbus_Mem_Alu_R[2]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1324z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1323z62958 (.O (px2966), .I0 (px3484), .I1 (p_nbus_Ex_D1[3]), .I2 (
         p_nbus_Mem_Alu_R[3]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1323z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1322z62958 (.O (px2967), .I0 (px3483), .I1 (p_nbus_Ex_D1[4]), .I2 (
         p_nbus_Mem_Alu_R[4]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1322z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1321z62958 (.O (px2968), .I0 (px3482), .I1 (p_nbus_Ex_D1[5]), .I2 (
         p_nbus_Mem_Alu_R[5]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1321z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1320z62958 (.O (px2969), .I0 (px3481), .I1 (p_nbus_Ex_D1[6]), .I2 (
         p_nbus_Mem_Alu_R[6]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1320z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1319z62958 (.O (px2970), .I0 (px3480), .I1 (p_nbus_Ex_D1[7]), .I2 (
         p_nbus_Mem_Alu_R[7]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1319z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1318z62958 (.O (px2971), .I0 (px3479), .I1 (p_nbus_Ex_D1[8]), .I2 (
         p_nbus_Mem_Alu_R[8]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1318z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1317z62958 (.O (px2972), .I0 (px3478), .I1 (p_nbus_Ex_D1[9]), .I2 (
         p_nbus_Mem_Alu_R[9]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (p_nbus_Ex_Fwd_A[1]
         )) ;
         defparam ix1317z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1316z62958 (.O (px2973), .I0 (px3477), .I1 (p_nbus_Ex_D1[10]), .I2 (
         p_nbus_Mem_Alu_R[10]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix1316z62958.INIT = 32'hCC55F0CC;
    LUT5 ix1315z62958 (.O (px2974), .I0 (px3476), .I1 (p_nbus_Ex_D1[11]), .I2 (
         p_nbus_Mem_Alu_R[11]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix1315z62958.INIT = 32'hCC55F0CC;
    LUT5 ix327z62958 (.O (px2975), .I0 (px3475), .I1 (p_nbus_Ex_D1[12]), .I2 (
         p_nbus_Mem_Alu_R[12]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix327z62958.INIT = 32'hCC55F0CC;
    LUT5 ix326z62958 (.O (px2976), .I0 (px3474), .I1 (p_nbus_Ex_D1[13]), .I2 (
         p_nbus_Mem_Alu_R[13]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix326z62958.INIT = 32'hCC55F0CC;
    LUT5 ix325z62958 (.O (px2977), .I0 (px3473), .I1 (p_nbus_Ex_D1[14]), .I2 (
         p_nbus_Mem_Alu_R[14]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix325z62958.INIT = 32'hCC55F0CC;
    LUT5 ix324z62958 (.O (px2978), .I0 (px3472), .I1 (p_nbus_Ex_D1[15]), .I2 (
         p_nbus_Mem_Alu_R[15]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix324z62958.INIT = 32'hCC55F0CC;
    LUT5 ix323z62958 (.O (px2979), .I0 (px3471), .I1 (p_nbus_Ex_D1[16]), .I2 (
         p_nbus_Mem_Alu_R[16]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix323z62958.INIT = 32'hCC55F0CC;
    LUT5 ix322z62958 (.O (px2980), .I0 (px3470), .I1 (p_nbus_Ex_D1[17]), .I2 (
         p_nbus_Mem_Alu_R[17]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix322z62958.INIT = 32'hCC55F0CC;
    LUT5 ix321z62958 (.O (px2981), .I0 (px3469), .I1 (p_nbus_Ex_D1[18]), .I2 (
         p_nbus_Mem_Alu_R[18]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix321z62958.INIT = 32'hCC55F0CC;
    LUT5 ix320z62958 (.O (px2982), .I0 (px3468), .I1 (p_nbus_Ex_D1[19]), .I2 (
         p_nbus_Mem_Alu_R[19]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix320z62958.INIT = 32'hCC55F0CC;
    LUT5 ix319z62958 (.O (px2983), .I0 (px3467), .I1 (p_nbus_Ex_D1[20]), .I2 (
         p_nbus_Mem_Alu_R[20]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix319z62958.INIT = 32'hCC55F0CC;
    LUT5 ix318z62958 (.O (px2984), .I0 (px3466), .I1 (p_nbus_Ex_D1[21]), .I2 (
         p_nbus_Mem_Alu_R[21]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix318z62958.INIT = 32'hCC55F0CC;
    LUT5 ix63490z62958 (.O (px2985), .I0 (px3465), .I1 (p_nbus_Ex_D1[22]), .I2 (
         p_nbus_Mem_Alu_R[22]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix63490z62958.INIT = 32'hCC55F0CC;
    LUT5 ix63491z62958 (.O (px2986), .I0 (px3464), .I1 (p_nbus_Ex_D1[23]), .I2 (
         p_nbus_Mem_Alu_R[23]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix63491z62958.INIT = 32'hCC55F0CC;
    LUT5 ix63492z62958 (.O (px2987), .I0 (px3463), .I1 (p_nbus_Ex_D1[24]), .I2 (
         p_nbus_Mem_Alu_R[24]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix63492z62958.INIT = 32'hCC55F0CC;
    LUT5 ix63493z62958 (.O (px2988), .I0 (px3462), .I1 (p_nbus_Ex_D1[25]), .I2 (
         p_nbus_Mem_Alu_R[25]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix63493z62958.INIT = 32'hCC55F0CC;
    LUT5 ix20409z62958 (.O (px2989), .I0 (nx20409z3), .I1 (p_nbus_Ex_D1[26]), .I2 (
         p_nbus_Mem_Alu_R[26]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix20409z62958.INIT = 32'hCC55F0CC;
    LUT5 ix20408z62958 (.O (px2990), .I0 (nx20408z3), .I1 (p_nbus_Ex_D1[27]), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix20408z62958.INIT = 32'hCC55F0CC;
    LUT5 ix20407z62958 (.O (px2991), .I0 (nx20407z3), .I1 (p_nbus_Ex_D1[28]), .I2 (
         p_nbus_Mem_Alu_R[28]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix20407z62958.INIT = 32'hCC55F0CC;
    LUT5 ix20406z62958 (.O (px2992), .I0 (nx20406z3), .I1 (p_nbus_Ex_D1[29]), .I2 (
         p_nbus_Mem_Alu_R[29]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix20406z62958.INIT = 32'hCC55F0CC;
    LUT5 ix20405z62958 (.O (px2993), .I0 (px3457), .I1 (p_nbus_Ex_D1[30]), .I2 (
         p_nbus_Mem_Alu_R[30]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix20405z62958.INIT = 32'hCC55F0CC;
    LUT6 ix20404z1313 (.O (px2994), .I0 (p_nbus_Wb_D[0]), .I1 (
         p_nbus_Wb_Alu_R[0]), .I2 (p_Wb_Reg2reg), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1]), .I5 (nx20404z3)) ;
         defparam ix20404z1313.INIT = 64'h00CA0000FFFFFFFF;
    LUT6 ix32963z2002 (.O (px3004), .I0 (px3288), .I1 (px3287), .I2 (px3436), .I3 (
         px3435), .I4 (nx32963z3), .I5 (alu_R_0n0s6[31])) ;
         defparam ix32963z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix32964z2002 (.O (px3005), .I0 (px3291), .I1 (px3290), .I2 (px3436), .I3 (
         px3435), .I4 (nx32964z3), .I5 (alu_R_0n0s6[30])) ;
         defparam ix32964z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix32965z2002 (.O (px3006), .I0 (px3294), .I1 (px3293), .I2 (px3436), .I3 (
         px3435), .I4 (nx32965z3), .I5 (alu_R_0n0s6[29])) ;
         defparam ix32965z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix32966z2002 (.O (px3007), .I0 (px3297), .I1 (px3296), .I2 (px3436), .I3 (
         px3435), .I4 (nx32966z3), .I5 (alu_R_0n0s6[28])) ;
         defparam ix32966z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix32967z2002 (.O (px3008), .I0 (px3300), .I1 (px3299), .I2 (px3436), .I3 (
         px3435), .I4 (nx32967z3), .I5 (alu_R_0n0s6[27])) ;
         defparam ix32967z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix32968z2002 (.O (px3009), .I0 (px3303), .I1 (px3302), .I2 (px3436), .I3 (
         px3435), .I4 (nx32968z3), .I5 (alu_R_0n0s6[26])) ;
         defparam ix32968z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33956z2002 (.O (px3010), .I0 (px3306), .I1 (px3305), .I2 (px3436), .I3 (
         px3435), .I4 (nx33956z3), .I5 (alu_R_0n0s6[25])) ;
         defparam ix33956z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33957z2002 (.O (px3011), .I0 (px3309), .I1 (px3308), .I2 (px3436), .I3 (
         px3435), .I4 (nx33957z3), .I5 (alu_R_0n0s6[24])) ;
         defparam ix33957z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33958z2002 (.O (px3012), .I0 (px3312), .I1 (px3311), .I2 (px3436), .I3 (
         px3435), .I4 (nx33958z3), .I5 (alu_R_0n0s6[23])) ;
         defparam ix33958z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33959z2002 (.O (px3013), .I0 (px3315), .I1 (px3314), .I2 (px3436), .I3 (
         px3435), .I4 (nx33959z3), .I5 (alu_R_0n0s6[22])) ;
         defparam ix33959z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33960z2002 (.O (px3014), .I0 (px3318), .I1 (px3317), .I2 (px3436), .I3 (
         px3435), .I4 (nx33960z3), .I5 (alu_R_0n0s6[21])) ;
         defparam ix33960z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33961z2002 (.O (px3015), .I0 (px3321), .I1 (px3320), .I2 (px3436), .I3 (
         px3435), .I4 (nx33961z3), .I5 (alu_R_0n0s6[20])) ;
         defparam ix33961z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33962z2002 (.O (px3016), .I0 (px3324), .I1 (px3323), .I2 (px3436), .I3 (
         px3435), .I4 (nx33962z3), .I5 (alu_R_0n0s6[19])) ;
         defparam ix33962z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33963z2002 (.O (px3017), .I0 (px3327), .I1 (px3326), .I2 (px3436), .I3 (
         px3435), .I4 (nx33963z3), .I5 (alu_R_0n0s6[18])) ;
         defparam ix33963z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33964z2002 (.O (px3018), .I0 (px3330), .I1 (px3329), .I2 (px3436), .I3 (
         px3435), .I4 (nx33964z3), .I5 (alu_R_0n0s6[17])) ;
         defparam ix33964z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix33965z2002 (.O (px3019), .I0 (px3333), .I1 (px3332), .I2 (px3436), .I3 (
         px3435), .I4 (nx33965z3), .I5 (alu_R_0n0s6[16])) ;
         defparam ix33965z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix34953z2002 (.O (px3020), .I0 (px3336), .I1 (px3335), .I2 (px3436), .I3 (
         px3435), .I4 (nx34953z3), .I5 (alu_R_0n0s6[15])) ;
         defparam ix34953z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix34954z2002 (.O (px3021), .I0 (px3339), .I1 (px3338), .I2 (px3436), .I3 (
         px3435), .I4 (nx34954z3), .I5 (alu_R_0n0s6[14])) ;
         defparam ix34954z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix34955z1682 (.O (px3022), .I0 (nx321z5), .I1 (px3341), .I2 (px3436), .I3 (
         px3435), .I4 (nx34955z3), .I5 (alu_R_0n0s6[13])) ;
         defparam ix34955z1682.INIT = 64'hFF7FF1700F7F0170;
    LUT6 ix34956z1682 (.O (px3023), .I0 (px3346), .I1 (px3345), .I2 (px3436), .I3 (
         px3435), .I4 (nx34956z3), .I5 (alu_R_0n0s6[12])) ;
         defparam ix34956z1682.INIT = 64'hF17FF170017F0170;
    LUT6 ix34957z1682 (.O (px3024), .I0 (px3350), .I1 (px3349), .I2 (px3436), .I3 (
         px3435), .I4 (nx34957z3), .I5 (alu_R_0n0s6[11])) ;
         defparam ix34957z1682.INIT = 64'hF17FF170017F0170;
    LUT6 ix34958z2002 (.O (px3025), .I0 (px3354), .I1 (px3353), .I2 (px3436), .I3 (
         px3435), .I4 (nx34958z3), .I5 (alu_R_0n0s6[10])) ;
         defparam ix34958z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix34959z2002 (.O (px3026), .I0 (px3357), .I1 (px3356), .I2 (px3436), .I3 (
         px3435), .I4 (nx34959z3), .I5 (alu_R_0n0s6[9])) ;
         defparam ix34959z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix34960z2002 (.O (px3027), .I0 (px3360), .I1 (px3359), .I2 (px3436), .I3 (
         px3435), .I4 (nx34960z3), .I5 (alu_R_0n0s6[8])) ;
         defparam ix34960z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix34961z2002 (.O (px3028), .I0 (px3363), .I1 (px3362), .I2 (px3436), .I3 (
         px3435), .I4 (nx34961z3), .I5 (alu_R_0n0s6[7])) ;
         defparam ix34961z2002.INIT = 64'hF2BFF2B002BF02B0;
    LUT6 ix34962z1682 (.O (px3029), .I0 (px3366), .I1 (px3365), .I2 (px3436), .I3 (
         px3435), .I4 (nx34962z3), .I5 (alu_R_0n0s6[1])) ;
         defparam ix34962z1682.INIT = 64'hF17FF170017F0170;
    LUT6 ix35950z1228 (.O (px3030), .I0 (nx35950z2), .I1 (px3369), .I2 (px3368)
         , .I3 (p_nbus_Ex_Aluc[0]), .I4 (p_nbus_Ex_Aluc[1]), .I5 (nx35950z5)) ;
         defparam ix35950z1228.INIT = 64'h00AE00AAFFAEFFAA;
    LUT6 ix35957z1682 (.O (px3037), .I0 (px3419), .I1 (nx35957z2), .I2 (px3436)
         , .I3 (px3435), .I4 (nx35957z3), .I5 (alu_R_0n0s6[2])) ;
         defparam ix35957z1682.INIT = 64'hF17FF170017F0170;
    LUT6 ix35958z1682 (.O (px3038), .I0 (px3423), .I1 (px3422), .I2 (px3436), .I3 (
         px3435), .I4 (nx35958z2), .I5 (alu_R_0n0s6[3])) ;
         defparam ix35958z1682.INIT = 64'hF17FF170017F0170;
    LUT6 ix35959z1682 (.O (px3039), .I0 (px3427), .I1 (px3426), .I2 (px3436), .I3 (
         px3435), .I4 (nx35959z2), .I5 (alu_R_0n0s6[4])) ;
         defparam ix35959z1682.INIT = 64'hF17FF170017F0170;
    LUT6 ix36947z1682 (.O (px3040), .I0 (px3431), .I1 (px3430), .I2 (px3436), .I3 (
         px3435), .I4 (nx36947z2), .I5 (alu_R_0n0s6[5])) ;
         defparam ix36947z1682.INIT = 64'hFF7FF1700F7F0170;
    LUT6 ix36948z1682 (.O (px3041), .I0 (nx36948z2), .I1 (nx36948z4), .I2 (
         px3436), .I3 (px3435), .I4 (nx36948z7), .I5 (alu_R_0n0s6[6])) ;
         defparam ix36948z1682.INIT = 64'hF17FF170017F0170;
    LUT4 ix60029z38200 (.O (nx60029z21), .I0 (px3419), .I1 (nx35957z2), .I2 (
         px3366), .I3 (px3365)) ;
         defparam ix60029z38200.INIT = 16'h9009;
    LUT6 ix60029z38199 (.O (nx60029z19), .I0 (nx36948z2), .I1 (nx36948z4), .I2 (
         px3346), .I3 (px3345), .I4 (nx321z5), .I5 (px3341)) ;
         defparam ix60029z38199.INIT = 64'h9009000000009009;
    LUT5 ix60029z1325 (.O (nx60029z18), .I0 (px3350), .I1 (px3349), .I2 (px3312)
         , .I3 (px3311), .I4 (nx63499z2)) ;
         defparam ix60029z1325.INIT = 32'h09900000;
    LUT6 ix14591z46316 (.O (nx14591z2), .I0 (p_nbus_Ex_D1[0]), .I1 (
         p_nbus_Mem_Alu_R[0]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3487), .I5 (px3288)) ;
         defparam ix14591z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix14590z46316 (.O (nx14590z2), .I0 (p_nbus_Ex_D1[1]), .I1 (
         p_nbus_Mem_Alu_R[1]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3486), .I5 (px3291)) ;
         defparam ix14590z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13602z46316 (.O (nx13602z2), .I0 (p_nbus_Ex_D1[2]), .I1 (
         p_nbus_Mem_Alu_R[2]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3485), .I5 (px3294)) ;
         defparam ix13602z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13601z46316 (.O (nx13601z2), .I0 (p_nbus_Ex_D1[3]), .I1 (
         p_nbus_Mem_Alu_R[3]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3484), .I5 (px3297)) ;
         defparam ix13601z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13600z46316 (.O (nx13600z2), .I0 (p_nbus_Ex_D1[4]), .I1 (
         p_nbus_Mem_Alu_R[4]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3483), .I5 (px3300)) ;
         defparam ix13600z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13599z46316 (.O (nx13599z2), .I0 (p_nbus_Ex_D1[5]), .I1 (
         p_nbus_Mem_Alu_R[5]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3482), .I5 (px3303)) ;
         defparam ix13599z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13598z46316 (.O (nx13598z2), .I0 (p_nbus_Ex_D1[6]), .I1 (
         p_nbus_Mem_Alu_R[6]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3481), .I5 (px3306)) ;
         defparam ix13598z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13597z46316 (.O (nx13597z2), .I0 (p_nbus_Ex_D1[7]), .I1 (
         p_nbus_Mem_Alu_R[7]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3480), .I5 (px3309)) ;
         defparam ix13597z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13596z46316 (.O (nx13596z2), .I0 (p_nbus_Ex_D1[8]), .I1 (
         p_nbus_Mem_Alu_R[8]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3479), .I5 (px3312)) ;
         defparam ix13596z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13595z46316 (.O (nx13595z2), .I0 (p_nbus_Ex_D1[9]), .I1 (
         p_nbus_Mem_Alu_R[9]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (p_nbus_Ex_Fwd_A[1]
         ), .I4 (px3478), .I5 (px3315)) ;
         defparam ix13595z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13594z46316 (.O (nx13594z2), .I0 (p_nbus_Ex_D1[10]), .I1 (
         p_nbus_Mem_Alu_R[10]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3477), .I5 (px3318)) ;
         defparam ix13594z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix13593z46316 (.O (nx13593z2), .I0 (p_nbus_Ex_D1[11]), .I1 (
         p_nbus_Mem_Alu_R[11]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3476), .I5 (px3321)) ;
         defparam ix13593z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix12605z46316 (.O (nx12605z2), .I0 (p_nbus_Ex_D1[12]), .I1 (
         p_nbus_Mem_Alu_R[12]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3475), .I5 (px3324)) ;
         defparam ix12605z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix12604z46316 (.O (nx12604z2), .I0 (p_nbus_Ex_D1[13]), .I1 (
         p_nbus_Mem_Alu_R[13]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3474), .I5 (px3327)) ;
         defparam ix12604z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix12603z46316 (.O (nx12603z2), .I0 (p_nbus_Ex_D1[14]), .I1 (
         p_nbus_Mem_Alu_R[14]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3473), .I5 (px3330)) ;
         defparam ix12603z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix12602z46316 (.O (nx12602z2), .I0 (p_nbus_Ex_D1[15]), .I1 (
         p_nbus_Mem_Alu_R[15]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3472), .I5 (px3333)) ;
         defparam ix12602z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix12601z46316 (.O (nx12601z2), .I0 (p_nbus_Ex_D1[16]), .I1 (
         p_nbus_Mem_Alu_R[16]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3471), .I5 (px3336)) ;
         defparam ix12601z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix12600z46316 (.O (nx12600z2), .I0 (p_nbus_Ex_D1[17]), .I1 (
         p_nbus_Mem_Alu_R[17]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3470), .I5 (px3339)) ;
         defparam ix12600z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix12599z21847 (.O (nx12599z2), .I0 (p_nbus_Ex_D1[18]), .I1 (
         p_nbus_Mem_Alu_R[18]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3469), .I5 (nx321z5)) ;
         defparam ix12599z21847.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix12598z21847 (.O (nx12598z2), .I0 (p_nbus_Ex_D1[19]), .I1 (
         p_nbus_Mem_Alu_R[19]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3468), .I5 (px3346)) ;
         defparam ix12598z21847.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix12597z21847 (.O (nx12597z2), .I0 (p_nbus_Ex_D1[20]), .I1 (
         p_nbus_Mem_Alu_R[20]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3467), .I5 (px3350)) ;
         defparam ix12597z21847.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix12596z46316 (.O (nx12596z2), .I0 (p_nbus_Ex_D1[21]), .I1 (
         p_nbus_Mem_Alu_R[21]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3466), .I5 (px3354)) ;
         defparam ix12596z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix39748z46316 (.O (nx39748z2), .I0 (p_nbus_Ex_D1[22]), .I1 (
         p_nbus_Mem_Alu_R[22]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3465), .I5 (px3357)) ;
         defparam ix39748z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix39749z46316 (.O (nx39749z2), .I0 (p_nbus_Ex_D1[23]), .I1 (
         p_nbus_Mem_Alu_R[23]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3464), .I5 (px3360)) ;
         defparam ix39749z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix39750z46316 (.O (nx39750z2), .I0 (p_nbus_Ex_D1[24]), .I1 (
         p_nbus_Mem_Alu_R[24]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3463), .I5 (px3363)) ;
         defparam ix39750z46316.INIT = 64'h5F355035A0CAAFCA;
    LUT6 ix39751z21847 (.O (nx39751z2), .I0 (p_nbus_Ex_D1[25]), .I1 (
         p_nbus_Mem_Alu_R[25]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3462), .I5 (nx36948z2)) ;
         defparam ix39751z21847.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix20409z21849 (.O (nx20409z4), .I0 (p_nbus_Ex_D1[26]), .I1 (
         p_nbus_Mem_Alu_R[26]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20409z3), .I5 (px3431)) ;
         defparam ix20409z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix20408z21849 (.O (nx20408z4), .I0 (p_nbus_Ex_D1[27]), .I1 (
         p_nbus_Mem_Alu_R[27]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20408z3), .I5 (px3427)) ;
         defparam ix20408z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix20407z21849 (.O (nx20407z4), .I0 (p_nbus_Ex_D1[28]), .I1 (
         p_nbus_Mem_Alu_R[28]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20407z3), .I5 (px3423)) ;
         defparam ix20407z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix20406z21849 (.O (nx20406z4), .I0 (p_nbus_Ex_D1[29]), .I1 (
         p_nbus_Mem_Alu_R[29]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (nx20406z3), .I5 (px3419)) ;
         defparam ix20406z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix20405z21849 (.O (nx20405z4), .I0 (p_nbus_Ex_D1[30]), .I1 (
         p_nbus_Mem_Alu_R[30]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1]), .I4 (px3457), .I5 (px3366)) ;
         defparam ix20405z21849.INIT = 64'hA0CAAFCA5F355035;
    LUT6 ix63499z10052 (.O (nx63499z2), .I0 (nx20404z3), .I1 (px3373), .I2 (
         px3371), .I3 (px3370), .I4 (\p_Ex_Extimm(0)  ), .I5 (p_Ex_Aluqb)) ;
         defparam ix63499z10052.INIT = 64'hDD2DDD2DDDDD2222;
    LUT2 ix32963z1319 (.O (nx32963z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[31])) ;
         defparam ix32963z1319.INIT = 4'h4;
    LUT6 ix2313z53541 (.O (px3288), .I0 (px3487), .I1 (p_nbus_Ex_D2[6]), .I2 (
         p_nbus_Mem_Alu_R[0]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix2313z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix32964z1319 (.O (nx32964z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[30])) ;
         defparam ix32964z1319.INIT = 4'h4;
    LUT6 ix2312z53541 (.O (px3291), .I0 (px3486), .I1 (p_nbus_Ex_D2[7]), .I2 (
         p_nbus_Mem_Alu_R[1]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix2312z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix32965z1319 (.O (nx32965z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[29])) ;
         defparam ix32965z1319.INIT = 4'h4;
    LUT6 ix1324z53541 (.O (px3294), .I0 (px3485), .I1 (p_nbus_Ex_D2[8]), .I2 (
         p_nbus_Mem_Alu_R[2]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1324z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix32966z1319 (.O (nx32966z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[28])) ;
         defparam ix32966z1319.INIT = 4'h4;
    LUT6 ix1323z53541 (.O (px3297), .I0 (px3484), .I1 (p_nbus_Ex_D2[9]), .I2 (
         p_nbus_Mem_Alu_R[3]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1323z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix32967z1319 (.O (nx32967z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[27])) ;
         defparam ix32967z1319.INIT = 4'h4;
    LUT6 ix1322z53541 (.O (px3300), .I0 (px3483), .I1 (p_nbus_Ex_D2[10]), .I2 (
         p_nbus_Mem_Alu_R[4]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1322z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix32968z1319 (.O (nx32968z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[26])) ;
         defparam ix32968z1319.INIT = 4'h4;
    LUT6 ix1321z53541 (.O (px3303), .I0 (px3482), .I1 (p_nbus_Ex_D2[11]), .I2 (
         p_nbus_Mem_Alu_R[5]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1321z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33956z1319 (.O (nx33956z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[25])) ;
         defparam ix33956z1319.INIT = 4'h4;
    LUT6 ix1320z53541 (.O (px3306), .I0 (px3481), .I1 (p_nbus_Ex_D2[12]), .I2 (
         p_nbus_Mem_Alu_R[6]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1320z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33957z1319 (.O (nx33957z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[24])) ;
         defparam ix33957z1319.INIT = 4'h4;
    LUT6 ix1319z53541 (.O (px3309), .I0 (px3480), .I1 (p_nbus_Ex_D2[13]), .I2 (
         p_nbus_Mem_Alu_R[7]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1319z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33958z1319 (.O (nx33958z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[23])) ;
         defparam ix33958z1319.INIT = 4'h4;
    LUT6 ix1318z53541 (.O (px3312), .I0 (px3479), .I1 (p_nbus_Ex_D2[14]), .I2 (
         p_nbus_Mem_Alu_R[8]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1318z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33959z1319 (.O (nx33959z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[22])) ;
         defparam ix33959z1319.INIT = 4'h4;
    LUT6 ix1317z53541 (.O (px3315), .I0 (px3478), .I1 (p_nbus_Ex_D2[15]), .I2 (
         p_nbus_Mem_Alu_R[9]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1317z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33960z1319 (.O (nx33960z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[21])) ;
         defparam ix33960z1319.INIT = 4'h4;
    LUT6 ix1316z53541 (.O (px3318), .I0 (px3477), .I1 (p_nbus_Ex_D2[16]), .I2 (
         p_nbus_Mem_Alu_R[10]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1316z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33961z1319 (.O (nx33961z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[20])) ;
         defparam ix33961z1319.INIT = 4'h4;
    LUT6 ix1315z53541 (.O (px3321), .I0 (px3476), .I1 (p_nbus_Ex_D2[17]), .I2 (
         p_nbus_Mem_Alu_R[11]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix1315z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33962z1319 (.O (nx33962z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[19])) ;
         defparam ix33962z1319.INIT = 4'h4;
    LUT6 ix327z53541 (.O (px3324), .I0 (px3475), .I1 (p_nbus_Ex_D2[18]), .I2 (
         p_nbus_Mem_Alu_R[12]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix327z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33963z1319 (.O (nx33963z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[18])) ;
         defparam ix33963z1319.INIT = 4'h4;
    LUT6 ix326z53541 (.O (px3327), .I0 (px3474), .I1 (p_nbus_Ex_D2[19]), .I2 (
         p_nbus_Mem_Alu_R[13]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix326z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33964z1319 (.O (nx33964z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[17])) ;
         defparam ix33964z1319.INIT = 4'h4;
    LUT6 ix325z53541 (.O (px3330), .I0 (px3473), .I1 (p_nbus_Ex_D2[20]), .I2 (
         p_nbus_Mem_Alu_R[14]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix325z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix33965z1319 (.O (nx33965z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[16])) ;
         defparam ix33965z1319.INIT = 4'h4;
    LUT6 ix324z53541 (.O (px3333), .I0 (px3472), .I1 (p_nbus_Ex_D2[21]), .I2 (
         p_nbus_Mem_Alu_R[15]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix324z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix34953z1319 (.O (nx34953z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[15])) ;
         defparam ix34953z1319.INIT = 4'h4;
    LUT6 ix323z53541 (.O (px3336), .I0 (px3471), .I1 (p_nbus_Ex_D2[22]), .I2 (
         p_nbus_Mem_Alu_R[16]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix323z53541.INIT = 64'hCC005500F000CC00;
    LUT2 ix34954z1319 (.O (nx34954z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[14])) ;
         defparam ix34954z1319.INIT = 4'h4;
    LUT6 ix322z53541 (.O (px3339), .I0 (px3470), .I1 (p_nbus_Ex_D2[23]), .I2 (
         p_nbus_Mem_Alu_R[17]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix322z53541.INIT = 64'hCC005500F000CC00;
    LUT3 ix34955z1331 (.O (nx34955z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         p_nbus_Ex_Aluc[1]), .I2 (alu_R_0n0s3[13])) ;
         defparam ix34955z1331.INIT = 8'h10;
    LUT6 ix321z44888 (.O (nx321z5), .I0 (px3343), .I1 (\p_Ex_Extimm(13)  ), .I2 (
         p_nbus_Mem_Alu_R[18]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix321z44888.INIT = 64'hAA33AA330A33AA33;
    LUT6 ix4321z23159 (.O (px3343), .I0 (p_nbus_Ex_D2[24]), .I1 (p_nbus_Wb_D[1])
         , .I2 (p_nbus_Wb_Alu_R[1]), .I3 (p_Wb_Reg2reg), .I4 (p_nbus_Ex_Fwd_B[0]
         ), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix4321z23159.INIT = 64'h55550F33FFFF5555;
    LUT2 ix34956z1319 (.O (nx34956z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[12])) ;
         defparam ix34956z1319.INIT = 4'h4;
    LUT2 ix34957z1319 (.O (nx34957z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[11])) ;
         defparam ix34957z1319.INIT = 4'h4;
    (* HLUTNM = "LUT62_4_1" *)
    LUT2 ix34958z1319 (.O (nx34958z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[10])) ;
         defparam ix34958z1319.INIT = 4'h4;
    LUT6 ix318z53541 (.O (px3354), .I0 (px3466), .I1 (p_nbus_Ex_D2[25]), .I2 (
         p_nbus_Mem_Alu_R[21]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix318z53541.INIT = 64'hCC005500F000CC00;
    (* HLUTNM = "LUT62_4_2" *)
    LUT2 ix34959z1319 (.O (nx34959z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[9])) ;
         defparam ix34959z1319.INIT = 4'h4;
    LUT6 ix63490z53541 (.O (px3357), .I0 (px3465), .I1 (p_nbus_Ex_D2[26]), .I2 (
         p_nbus_Mem_Alu_R[22]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix63490z53541.INIT = 64'hCC005500F000CC00;
    (* HLUTNM = "LUT62_4_2" *)
    LUT2 ix34960z1319 (.O (nx34960z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[8])) ;
         defparam ix34960z1319.INIT = 4'h4;
    LUT6 ix63491z53541 (.O (px3360), .I0 (px3464), .I1 (p_nbus_Ex_D2[27]), .I2 (
         p_nbus_Mem_Alu_R[23]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix63491z53541.INIT = 64'hCC005500F000CC00;
    (* HLUTNM = "LUT62_4_3" *)
    LUT2 ix34961z1319 (.O (nx34961z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[7])) ;
         defparam ix34961z1319.INIT = 4'h4;
    LUT6 ix63492z53541 (.O (px3363), .I0 (px3463), .I1 (p_nbus_Ex_D2[28]), .I2 (
         p_nbus_Mem_Alu_R[24]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix63492z53541.INIT = 64'hCC005500F000CC00;
    (* HLUTNM = "LUT62_4_3" *)
    LUT2 ix34962z1319 (.O (nx34962z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[1])) ;
         defparam ix34962z1319.INIT = 4'h4;
    LUT5 ix20404z1319 (.O (px3370), .I0 (p_nbus_Wb_D[0]), .I1 (
         p_nbus_Wb_Alu_R[0]), .I2 (p_Wb_Reg2reg), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix20404z1319.INIT = 32'h00CA0000;
    LUT4 ix20404z25691 (.O (px3371), .I0 (p_nbus_Ex_D2[29]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (p_nbus_Ex_Fwd_B[0]), .I3 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix20404z25691.INIT = 16'h5F35;
    LUT6 ix35950z54563 (.O (nx35950z2), .I0 (nx20404z3), .I1 (px3373), .I2 (
         p_nbus_Ex_Aluc[1]), .I3 (p_nbus_Ex_Aluc[2]), .I4 (alu_R_0n0s3[0]), .I5 (
         alu_R_0n0s6[0])) ;
         defparam ix35950z54563.INIT = 64'hDF0FDF00D00FD000;
    LUT5 ix20404z1317 (.O (px3373), .I0 (p_nbus_Wb_D[0]), .I1 (
         p_nbus_Wb_Alu_R[0]), .I2 (p_Wb_Reg2reg), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix20404z1317.INIT = 32'h00CA0000;
    LUT4 ix20404z25688 (.O (nx20404z3), .I0 (p_nbus_Ex_D1[31]), .I1 (
         p_nbus_Mem_Alu_R[31]), .I2 (p_nbus_Ex_Fwd_A[0]), .I3 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix20404z25688.INIT = 16'h5F35;
    (* HLUTNM = "LUT62_4_4" *)
    LUT2 ix35957z1320 (.O (nx35957z3), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[2])) ;
         defparam ix35957z1320.INIT = 4'h4;
    LUT5 ix35957z5206 (.O (nx35957z2), .I0 (nx20406z3), .I1 (p_nbus_Ex_D1[29]), 
         .I2 (p_nbus_Mem_Alu_R[29]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix35957z5206.INIT = 32'h33AA0F33;
    LUT6 ix13293z1313 (.O (px3420), .I0 (p_nbus_Mem_Alu_R[29]), .I1 (
         p_nbus_Wb_D[2]), .I2 (p_nbus_Wb_Alu_R[2]), .I3 (p_Wb_Reg2reg), .I4 (
         p_nbus_Ex_Fwd_B[0]), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix13293z1313.INIT = 64'hFFFF0F335555FFFF;
    (* HLUTNM = "LUT62_4_4" *)
    LUT2 ix35958z1319 (.O (nx35958z2), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[3])) ;
         defparam ix35958z1319.INIT = 4'h4;
    LUT5 ix13295z5205 (.O (px3422), .I0 (nx20407z3), .I1 (p_nbus_Ex_D1[28]), .I2 (
         p_nbus_Mem_Alu_R[28]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix13295z5205.INIT = 32'h33AA0F33;
    LUT6 ix13297z1313 (.O (px3424), .I0 (p_nbus_Mem_Alu_R[28]), .I1 (
         p_nbus_Wb_D[3]), .I2 (p_nbus_Wb_Alu_R[3]), .I3 (p_Wb_Reg2reg), .I4 (
         p_nbus_Ex_Fwd_B[0]), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix13297z1313.INIT = 64'hFFFF0F335555FFFF;
    (* HLUTNM = "LUT62_4_5" *)
    LUT2 ix35959z1319 (.O (nx35959z2), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[4])) ;
         defparam ix35959z1319.INIT = 4'h4;
    LUT5 ix13299z5205 (.O (px3426), .I0 (nx20408z3), .I1 (p_nbus_Ex_D1[27]), .I2 (
         p_nbus_Mem_Alu_R[27]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix13299z5205.INIT = 32'h33AA0F33;
    LUT6 ix13301z1313 (.O (px3428), .I0 (p_nbus_Mem_Alu_R[27]), .I1 (
         p_nbus_Wb_D[4]), .I2 (p_nbus_Wb_Alu_R[4]), .I3 (p_Wb_Reg2reg), .I4 (
         p_nbus_Ex_Fwd_B[0]), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix13301z1313.INIT = 64'hFFFF0F335555FFFF;
    (* HLUTNM = "LUT62_4_1" *)
    LUT3 ix36947z1331 (.O (nx36947z2), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         p_nbus_Ex_Aluc[1]), .I2 (alu_R_0n0s3[5])) ;
         defparam ix36947z1331.INIT = 8'h10;
    LUT5 ix14290z5205 (.O (px3430), .I0 (nx20409z3), .I1 (p_nbus_Ex_D1[26]), .I2 (
         p_nbus_Mem_Alu_R[26]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix14290z5205.INIT = 32'h33AA0F33;
    LUT6 ix20409z44888 (.O (px3431), .I0 (px3432), .I1 (\p_Ex_Extimm(13)  ), .I2 (
         p_nbus_Mem_Alu_R[26]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix20409z44888.INIT = 64'hAA33AA330A33AA33;
    LUT6 ix14292z23159 (.O (px3432), .I0 (p_nbus_Ex_D2[30]), .I1 (p_nbus_Wb_D[5]
         ), .I2 (p_nbus_Wb_Alu_R[5]), .I3 (p_Wb_Reg2reg), .I4 (
         p_nbus_Ex_Fwd_B[0]), .I5 (p_nbus_Ex_Fwd_B[1])) ;
         defparam ix14292z23159.INIT = 64'h55550F33FFFF5555;
    (* HLUTNM = "LUT62_4_5" *)
    LUT2 ix36948z1322 (.O (nx36948z7), .I0 (p_nbus_Ex_Aluc[0]), .I1 (
         alu_R_0n0s3[6])) ;
         defparam ix36948z1322.INIT = 4'h4;
    LUT5 ix36948z5208 (.O (nx36948z4), .I0 (px3462), .I1 (p_nbus_Ex_D1[25]), .I2 (
         p_nbus_Mem_Alu_R[25]), .I3 (p_nbus_Ex_Fwd_A[0]), .I4 (
         p_nbus_Ex_Fwd_A[1])) ;
         defparam ix36948z5208.INIT = 32'h33AA0F33;
    LUT6 ix36948z53554 (.O (nx36948z2), .I0 (px3462), .I1 (px3439), .I2 (
         \p_Ex_Op(0)  ), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix36948z53554.INIT = 64'hCC0F880FCC0FCC0F;
    LUT4 ix14299z25687 (.O (px3439), .I0 (p_nbus_Ex_D2[31]), .I1 (
         p_nbus_Mem_Alu_R[25]), .I2 (p_nbus_Ex_Fwd_B[0]), .I3 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix14299z25687.INIT = 16'h5F35;
    LUT3 ix20405z1368 (.O (px3457), .I0 (p_nbus_Wb_D[6]), .I1 (
         p_nbus_Wb_Alu_R[6]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix20405z1368.INIT = 8'h35;
    LUT3 ix20406z1368 (.O (nx20406z3), .I0 (p_nbus_Wb_D[2]), .I1 (
         p_nbus_Wb_Alu_R[2]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix20406z1368.INIT = 8'h35;
    LUT3 ix20407z1368 (.O (nx20407z3), .I0 (p_nbus_Wb_D[3]), .I1 (
         p_nbus_Wb_Alu_R[3]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix20407z1368.INIT = 8'h35;
    LUT3 ix20408z1368 (.O (nx20408z3), .I0 (p_nbus_Wb_D[4]), .I1 (
         p_nbus_Wb_Alu_R[4]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix20408z1368.INIT = 8'h35;
    LUT3 ix20409z1368 (.O (nx20409z3), .I0 (p_nbus_Wb_D[5]), .I1 (
         p_nbus_Wb_Alu_R[5]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix20409z1368.INIT = 8'h35;
    LUT3 ix36948z1369 (.O (px3462), .I0 (p_nbus_Wb_D[7]), .I1 (
         p_nbus_Wb_Alu_R[7]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix36948z1369.INIT = 8'h35;
    LUT3 ix63492z1368 (.O (px3463), .I0 (p_nbus_Wb_D[8]), .I1 (
         p_nbus_Wb_Alu_R[8]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix63492z1368.INIT = 8'h35;
    LUT3 ix63491z1368 (.O (px3464), .I0 (p_nbus_Wb_D[9]), .I1 (
         p_nbus_Wb_Alu_R[9]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix63491z1368.INIT = 8'h35;
    LUT3 ix63490z1368 (.O (px3465), .I0 (p_nbus_Wb_D[10]), .I1 (
         p_nbus_Wb_Alu_R[10]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix63490z1368.INIT = 8'h35;
    LUT3 ix318z1368 (.O (px3466), .I0 (p_nbus_Wb_D[11]), .I1 (
         p_nbus_Wb_Alu_R[11]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix318z1368.INIT = 8'h35;
    LUT3 ix319z1368 (.O (px3467), .I0 (p_nbus_Wb_D[12]), .I1 (
         p_nbus_Wb_Alu_R[12]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix319z1368.INIT = 8'h35;
    LUT3 ix320z1368 (.O (px3468), .I0 (p_nbus_Wb_D[13]), .I1 (
         p_nbus_Wb_Alu_R[13]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix320z1368.INIT = 8'h35;
    LUT3 ix321z1368 (.O (px3469), .I0 (p_nbus_Wb_D[1]), .I1 (p_nbus_Wb_Alu_R[1])
         , .I2 (p_Wb_Reg2reg)) ;
         defparam ix321z1368.INIT = 8'h35;
    LUT3 ix322z1368 (.O (px3470), .I0 (p_nbus_Wb_D[14]), .I1 (
         p_nbus_Wb_Alu_R[14]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix322z1368.INIT = 8'h35;
    LUT3 ix323z1368 (.O (px3471), .I0 (p_nbus_Wb_D[15]), .I1 (
         p_nbus_Wb_Alu_R[15]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix323z1368.INIT = 8'h35;
    LUT3 ix324z1368 (.O (px3472), .I0 (p_nbus_Wb_D[16]), .I1 (
         p_nbus_Wb_Alu_R[16]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix324z1368.INIT = 8'h35;
    LUT3 ix325z1368 (.O (px3473), .I0 (p_nbus_Wb_D[17]), .I1 (
         p_nbus_Wb_Alu_R[17]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix325z1368.INIT = 8'h35;
    LUT3 ix326z1368 (.O (px3474), .I0 (p_nbus_Wb_D[18]), .I1 (
         p_nbus_Wb_Alu_R[18]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix326z1368.INIT = 8'h35;
    LUT3 ix327z1368 (.O (px3475), .I0 (p_nbus_Wb_D[19]), .I1 (
         p_nbus_Wb_Alu_R[19]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix327z1368.INIT = 8'h35;
    LUT3 ix1315z1368 (.O (px3476), .I0 (p_nbus_Wb_D[20]), .I1 (
         p_nbus_Wb_Alu_R[20]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1315z1368.INIT = 8'h35;
    LUT3 ix1316z1368 (.O (px3477), .I0 (p_nbus_Wb_D[21]), .I1 (
         p_nbus_Wb_Alu_R[21]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1316z1368.INIT = 8'h35;
    LUT3 ix1317z1368 (.O (px3478), .I0 (p_nbus_Wb_D[22]), .I1 (
         p_nbus_Wb_Alu_R[22]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1317z1368.INIT = 8'h35;
    LUT3 ix1318z1368 (.O (px3479), .I0 (p_nbus_Wb_D[23]), .I1 (
         p_nbus_Wb_Alu_R[23]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1318z1368.INIT = 8'h35;
    LUT3 ix1319z1368 (.O (px3480), .I0 (p_nbus_Wb_D[24]), .I1 (
         p_nbus_Wb_Alu_R[24]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1319z1368.INIT = 8'h35;
    LUT3 ix1320z1368 (.O (px3481), .I0 (p_nbus_Wb_D[25]), .I1 (
         p_nbus_Wb_Alu_R[25]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1320z1368.INIT = 8'h35;
    LUT3 ix1321z1368 (.O (px3482), .I0 (p_nbus_Wb_D[26]), .I1 (
         p_nbus_Wb_Alu_R[26]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1321z1368.INIT = 8'h35;
    LUT3 ix1322z1368 (.O (px3483), .I0 (p_nbus_Wb_D[27]), .I1 (
         p_nbus_Wb_Alu_R[27]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1322z1368.INIT = 8'h35;
    LUT3 ix1323z1368 (.O (px3484), .I0 (p_nbus_Wb_D[28]), .I1 (
         p_nbus_Wb_Alu_R[28]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1323z1368.INIT = 8'h35;
    LUT3 ix1324z1368 (.O (px3485), .I0 (p_nbus_Wb_D[29]), .I1 (
         p_nbus_Wb_Alu_R[29]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix1324z1368.INIT = 8'h35;
    LUT3 ix2312z1368 (.O (px3486), .I0 (p_nbus_Wb_D[30]), .I1 (
         p_nbus_Wb_Alu_R[30]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix2312z1368.INIT = 8'h35;
    LUT3 ix2313z1368 (.O (px3487), .I0 (p_nbus_Wb_D[31]), .I1 (
         p_nbus_Wb_Alu_R[31]), .I2 (p_Wb_Reg2reg)) ;
         defparam ix2313z1368.INIT = 8'h35;
    MUXCY R_add32_0i1_muxcy_0 (.O (nx20405z1), .CI (px2857), .DI (px2994), .S (
          nx20404z4)) ;
    MUXCY R_add32_0i1_muxcy_1 (.O (nx20406z1), .CI (nx20405z1), .DI (px2993), .S (
          nx20405z4)) ;
    MUXCY R_add32_0i1_muxcy_2 (.O (nx20407z1), .CI (nx20406z1), .DI (px2992), .S (
          nx20406z4)) ;
    MUXCY R_add32_0i1_muxcy_3 (.O (nx20408z1), .CI (nx20407z1), .DI (px2991), .S (
          nx20407z4)) ;
    MUXCY R_add32_0i1_muxcy_4 (.O (nx20409z1), .CI (nx20408z1), .DI (px2990), .S (
          nx20408z4)) ;
    MUXCY R_add32_0i1_muxcy_5 (.O (nx39751z1), .CI (nx20409z1), .DI (px2989), .S (
          nx20409z4)) ;
    MUXCY R_add32_0i1_muxcy_6 (.O (nx39750z1), .CI (nx39751z1), .DI (px2988), .S (
          nx39751z2)) ;
    MUXCY R_add32_0i1_muxcy_7 (.O (nx39749z1), .CI (nx39750z1), .DI (px2987), .S (
          nx39750z2)) ;
    MUXCY R_add32_0i1_muxcy_8 (.O (nx39748z1), .CI (nx39749z1), .DI (px2986), .S (
          nx39749z2)) ;
    MUXCY R_add32_0i1_muxcy_9 (.O (nx12596z1), .CI (nx39748z1), .DI (px2985), .S (
          nx39748z2)) ;
    MUXCY R_add32_0i1_muxcy_10 (.O (nx12597z1), .CI (nx12596z1), .DI (px2984), .S (
          nx12596z2)) ;
    MUXCY R_add32_0i1_muxcy_11 (.O (nx12598z1), .CI (nx12597z1), .DI (px2983), .S (
          nx12597z2)) ;
    MUXCY R_add32_0i1_muxcy_12 (.O (nx12599z1), .CI (nx12598z1), .DI (px2982), .S (
          nx12598z2)) ;
    MUXCY R_add32_0i1_muxcy_13 (.O (nx12600z1), .CI (nx12599z1), .DI (px2981), .S (
          nx12599z2)) ;
    MUXCY R_add32_0i1_muxcy_14 (.O (nx12601z1), .CI (nx12600z1), .DI (px2980), .S (
          nx12600z2)) ;
    MUXCY R_add32_0i1_muxcy_15 (.O (nx12602z1), .CI (nx12601z1), .DI (px2979), .S (
          nx12601z2)) ;
    MUXCY R_add32_0i1_muxcy_16 (.O (nx12603z1), .CI (nx12602z1), .DI (px2978), .S (
          nx12602z2)) ;
    MUXCY R_add32_0i1_muxcy_17 (.O (nx12604z1), .CI (nx12603z1), .DI (px2977), .S (
          nx12603z2)) ;
    MUXCY R_add32_0i1_muxcy_18 (.O (nx12605z1), .CI (nx12604z1), .DI (px2976), .S (
          nx12604z2)) ;
    MUXCY R_add32_0i1_muxcy_19 (.O (nx13593z1), .CI (nx12605z1), .DI (px2975), .S (
          nx12605z2)) ;
    MUXCY R_add32_0i1_muxcy_20 (.O (nx13594z1), .CI (nx13593z1), .DI (px2974), .S (
          nx13593z2)) ;
    MUXCY R_add32_0i1_muxcy_21 (.O (nx13595z1), .CI (nx13594z1), .DI (px2973), .S (
          nx13594z2)) ;
    MUXCY R_add32_0i1_muxcy_22 (.O (nx13596z1), .CI (nx13595z1), .DI (px2972), .S (
          nx13595z2)) ;
    MUXCY R_add32_0i1_muxcy_23 (.O (nx13597z1), .CI (nx13596z1), .DI (px2971), .S (
          nx13596z2)) ;
    MUXCY R_add32_0i1_muxcy_24 (.O (nx13598z1), .CI (nx13597z1), .DI (px2970), .S (
          nx13597z2)) ;
    MUXCY R_add32_0i1_muxcy_25 (.O (nx13599z1), .CI (nx13598z1), .DI (px2969), .S (
          nx13598z2)) ;
    MUXCY R_add32_0i1_muxcy_26 (.O (nx13600z1), .CI (nx13599z1), .DI (px2968), .S (
          nx13599z2)) ;
    MUXCY R_add32_0i1_muxcy_27 (.O (nx13601z1), .CI (nx13600z1), .DI (px2967), .S (
          nx13600z2)) ;
    MUXCY R_add32_0i1_muxcy_28 (.O (nx13602z1), .CI (nx13601z1), .DI (px2966), .S (
          nx13601z2)) ;
    MUXCY R_add32_0i1_muxcy_29 (.O (nx14590z1), .CI (nx13602z1), .DI (px2965), .S (
          nx13602z2)) ;
    MUXCY R_add32_0i1_muxcy_30 (.O (nx14591z1), .CI (nx14590z1), .DI (px2964), .S (
          nx14590z2)) ;
    MUXCY Z_eq_0_ix60029z63350 (.O (nx60029z10), .CI (px2855), .DI (px2857), .S (
          px3215)) ;
    MUXCY Z_eq_0_ix60029z63349 (.O (nx60029z9), .CI (nx60029z10), .DI (px2857), 
          .S (px3214)) ;
    MUXCY Z_eq_0_ix60029z63348 (.O (nx60029z8), .CI (nx60029z9), .DI (px2857), .S (
          px3213)) ;
    MUXCY Z_eq_0_ix60029z63347 (.O (nx60029z7), .CI (nx60029z8), .DI (px2857), .S (
          px3212)) ;
    MUXCY Z_eq_0_ix60029z63346 (.O (nx60029z6), .CI (nx60029z7), .DI (px2857), .S (
          px3211)) ;
    MUXCY Z_eq_0_ix60029z63345 (.O (nx60029z5), .CI (nx60029z6), .DI (px2857), .S (
          px3210)) ;
    MUXCY Z_eq_0_ix60029z63344 (.O (nx60029z4), .CI (nx60029z5), .DI (px2857), .S (
          px3209)) ;
    MUXCY Z_eq_0_ix60029z63343 (.O (nx60029z3), .CI (nx60029z4), .DI (px2857), .S (
          nx60029z18)) ;
    MUXCY Z_eq_0_ix60029z63342 (.O (nx60029z2), .CI (nx60029z3), .DI (px2857), .S (
          nx60029z19)) ;
    MUXCY Z_eq_0_ix60029z63341 (.O (nx60029z1), .CI (nx60029z2), .DI (px2857), .S (
          px3206)) ;
    MUXCY R_sub32_0i5_muxcy_0 (.O (nx63498z1), .CI (px2855), .DI (px2994), .S (
          nx63499z2)) ;
    MUXCY R_sub32_0i5_muxcy_1 (.O (nx63497z1), .CI (nx63498z1), .DI (px2993), .S (
          nx63498z2)) ;
    MUXCY R_sub32_0i5_muxcy_2 (.O (nx63496z1), .CI (nx63497z1), .DI (px2992), .S (
          nx63497z2)) ;
    MUXCY R_sub32_0i5_muxcy_3 (.O (nx63495z1), .CI (nx63496z1), .DI (px2991), .S (
          nx63496z2)) ;
    MUXCY R_sub32_0i5_muxcy_4 (.O (nx63494z1), .CI (nx63495z1), .DI (px2990), .S (
          nx63495z2)) ;
    MUXCY R_sub32_0i5_muxcy_5 (.O (nx58118z1), .CI (nx63494z1), .DI (px2989), .S (
          nx63494z2)) ;
    MUXCY R_sub32_0i5_muxcy_6 (.O (nx63492z1), .CI (nx58118z1), .DI (px2988), .S (
          nx58118z2)) ;
    MUXCY R_sub32_0i5_muxcy_7 (.O (nx63491z1), .CI (nx63492z1), .DI (px2987), .S (
          nx63492z4)) ;
    MUXCY R_sub32_0i5_muxcy_8 (.O (nx63490z1), .CI (nx63491z1), .DI (px2986), .S (
          nx63491z4)) ;
    MUXCY R_sub32_0i5_muxcy_9 (.O (nx318z1), .CI (nx63490z1), .DI (px2985), .S (
          nx63490z4)) ;
    MUXCY R_sub32_0i5_muxcy_10 (.O (nx319z1), .CI (nx318z1), .DI (px2984), .S (
          nx318z4)) ;
    MUXCY R_sub32_0i5_muxcy_11 (.O (nx320z1), .CI (nx319z1), .DI (px2983), .S (
          nx319z4)) ;
    MUXCY R_sub32_0i5_muxcy_12 (.O (nx321z1), .CI (nx320z1), .DI (px2982), .S (
          nx320z4)) ;
    MUXCY R_sub32_0i5_muxcy_13 (.O (nx322z1), .CI (nx321z1), .DI (px2981), .S (
          nx321z4)) ;
    MUXCY R_sub32_0i5_muxcy_14 (.O (nx323z1), .CI (nx322z1), .DI (px2980), .S (
          nx322z4)) ;
    MUXCY R_sub32_0i5_muxcy_15 (.O (nx324z1), .CI (nx323z1), .DI (px2979), .S (
          nx323z4)) ;
    MUXCY R_sub32_0i5_muxcy_16 (.O (nx325z1), .CI (nx324z1), .DI (px2978), .S (
          nx324z4)) ;
    MUXCY R_sub32_0i5_muxcy_17 (.O (nx326z1), .CI (nx325z1), .DI (px2977), .S (
          nx325z4)) ;
    MUXCY R_sub32_0i5_muxcy_18 (.O (nx327z1), .CI (nx326z1), .DI (px2976), .S (
          nx326z4)) ;
    MUXCY R_sub32_0i5_muxcy_19 (.O (nx1315z1), .CI (nx327z1), .DI (px2975), .S (
          nx327z4)) ;
    MUXCY R_sub32_0i5_muxcy_20 (.O (nx1316z1), .CI (nx1315z1), .DI (px2974), .S (
          nx1315z4)) ;
    MUXCY R_sub32_0i5_muxcy_21 (.O (nx1317z1), .CI (nx1316z1), .DI (px2973), .S (
          nx1316z4)) ;
    MUXCY R_sub32_0i5_muxcy_22 (.O (nx1318z1), .CI (nx1317z1), .DI (px2972), .S (
          nx1317z4)) ;
    MUXCY R_sub32_0i5_muxcy_23 (.O (nx1319z1), .CI (nx1318z1), .DI (px2971), .S (
          nx1318z4)) ;
    MUXCY R_sub32_0i5_muxcy_24 (.O (nx1320z1), .CI (nx1319z1), .DI (px2970), .S (
          nx1319z4)) ;
    MUXCY R_sub32_0i5_muxcy_25 (.O (nx1321z1), .CI (nx1320z1), .DI (px2969), .S (
          nx1320z4)) ;
    MUXCY R_sub32_0i5_muxcy_26 (.O (nx1322z1), .CI (nx1321z1), .DI (px2968), .S (
          nx1321z4)) ;
    MUXCY R_sub32_0i5_muxcy_27 (.O (nx1323z1), .CI (nx1322z1), .DI (px2967), .S (
          nx1322z4)) ;
    MUXCY R_sub32_0i5_muxcy_28 (.O (nx1324z1), .CI (nx1323z1), .DI (px2966), .S (
          nx1323z4)) ;
    MUXCY R_sub32_0i5_muxcy_29 (.O (nx2312z1), .CI (nx1324z1), .DI (px2965), .S (
          nx1324z4)) ;
    MUXCY R_sub32_0i5_muxcy_30 (.O (nx2313z1), .CI (nx2312z1), .DI (px2964), .S (
          nx2312z4)) ;
endmodule


module ID_EX_unfolded0_0 ( \p_Rs_1_0(0)  , \p_Rs_1_0(1)  , \p_Rs_1_0(2)  , 
                           px3449, p_CLR_N_int, px3450, px3452, px3419, px3370, 
                           px3371, px3369, px3366, px3350, px3346, px3422, 
                           px3423, px3426, px3427, px3430, px3431, px3206, 
                           px3367, p_nbus_Ex_D2, px3003, px3420, px3002, px3424, 
                           px3001, px3428, px3000, p_nbus_Mem_Alu_R, px3432, 
                           px2999, px3439, px3462, px2998, px3351, px2997, 
                           px3347, px2996, px3343, px2995, \p_Pc_Add4(31)  , 
                           px2962, \p_Pc_Add4(30)  , px2960, \p_Pc_Add4(29)  , 
                           px2958, \p_Pc_Add4(28)  , px2956, \p_Pc_Add4(27)  , 
                           px2954, \p_Pc_Add4(26)  , px2952, \p_Pc_Add4(25)  , 
                           px2950, \p_Pc_Add4(24)  , px2948, \p_Pc_Add4(23)  , 
                           px2946, \p_Pc_Add4(22)  , px2944, \p_Pc_Add4(21)  , 
                           px2942, \p_Pc_Add4(20)  , px2940, \p_Pc_Add4(19)  , 
                           px2938, \p_Pc_Add4(18)  , px2936, \p_Pc_Add4(17)  , 
                           px2934, \p_Pc_Add4(16)  , px2932, \p_Pc_Add4(15)  , 
                           px2930, \p_Pc_Add4(14)  , px2928, \p_Pc_Add4(13)  , 
                           px2926, \p_Pc_Add4(12)  , px2924, \p_Pc_Add4(11)  , 
                           px2922, \p_Pc_Add4(10)  , px2920, \p_Pc_Add4(9)  , 
                           px2918, \p_Pc_Add4(8)  , px2916, \p_Pc_Add4(7)  , 
                           px2914, \p_Pc_Add4(6)  , px2912, \p_Pc_Add4(5)  , 
                           px2910, \p_Pc_Add4(4)  , px2908, \p_Pc_Add4(3)  , 
                           px2906, \p_Pc_Add4(2)  , px2904, p_nbus_Addr_1_0, 
                           px2902, p_Ex_Z, px2900, \p_Rt_1_0(2)  , \p_Rt_1_0(1)  , 
                           \p_Rt_1_0(0)  , \p_Id_Extimm(0)  , \p_Ex_Extimm(0)  , 
                           \p_Id_Extimm(1)  , \p_Id_Extimm(2)  , 
                           \p_Id_Extimm(3)  , \p_Id_Extimm(4)  , 
                           \p_Id_Extimm(13)  , \p_Ex_Extimm(13)  , 
                           \p_Id_Inst(26)  , \p_Ex_Op(0)  , \p_Id_Extimm(11)  , 
                           \p_Id_Extimm(12)  , \p_Id_Inst(28)  , \p_Id_Inst(29)  , 
                           p_nbus_Ex_Rd, p_nbus_Ex_Aluc, px3253, p_nbus_Ex_Fwd_A, 
                           px3255, px3256, p_nbus_Ex_Fwd_B, px3258, p_Ex_Wreg, 
                           p_Ex_Reg2reg, p_Ex_Wmem, p_Ex_Aluqb, 
                           p_nbus_Id_Pc_Add4, px3444, p_EN_int, p_CLK_int, 
                           px2857 ) ;

    input \p_Rs_1_0(0)   ;
    input \p_Rs_1_0(1)   ;
    input \p_Rs_1_0(2)   ;
    output px3449 ;
    input p_CLR_N_int ;
    output px3450 ;
    output px3452 ;
    output px3419 ;
    input px3370 ;
    input px3371 ;
    output px3369 ;
    output px3366 ;
    output px3350 ;
    output px3346 ;
    input px3422 ;
    output px3423 ;
    input px3426 ;
    output px3427 ;
    input px3430 ;
    input px3431 ;
    output px3206 ;
    input px3367 ;
    input [31:26]p_nbus_Ex_D2 ;
    output px3003 ;
    input px3420 ;
    output px3002 ;
    input px3424 ;
    output px3001 ;
    input px3428 ;
    output px3000 ;
    input [31:30]p_nbus_Mem_Alu_R ;
    input px3432 ;
    output px2999 ;
    input px3439 ;
    input px3462 ;
    output px2998 ;
    input px3351 ;
    output px2997 ;
    input px3347 ;
    output px2996 ;
    input px3343 ;
    output px2995 ;
    input \p_Pc_Add4(31)   ;
    output px2962 ;
    input \p_Pc_Add4(30)   ;
    output px2960 ;
    input \p_Pc_Add4(29)   ;
    output px2958 ;
    input \p_Pc_Add4(28)   ;
    output px2956 ;
    input \p_Pc_Add4(27)   ;
    output px2954 ;
    input \p_Pc_Add4(26)   ;
    output px2952 ;
    input \p_Pc_Add4(25)   ;
    output px2950 ;
    input \p_Pc_Add4(24)   ;
    output px2948 ;
    input \p_Pc_Add4(23)   ;
    output px2946 ;
    input \p_Pc_Add4(22)   ;
    output px2944 ;
    input \p_Pc_Add4(21)   ;
    output px2942 ;
    input \p_Pc_Add4(20)   ;
    output px2940 ;
    input \p_Pc_Add4(19)   ;
    output px2938 ;
    input \p_Pc_Add4(18)   ;
    output px2936 ;
    input \p_Pc_Add4(17)   ;
    output px2934 ;
    input \p_Pc_Add4(16)   ;
    output px2932 ;
    input \p_Pc_Add4(15)   ;
    output px2930 ;
    input \p_Pc_Add4(14)   ;
    output px2928 ;
    input \p_Pc_Add4(13)   ;
    output px2926 ;
    input \p_Pc_Add4(12)   ;
    output px2924 ;
    input \p_Pc_Add4(11)   ;
    output px2922 ;
    input \p_Pc_Add4(10)   ;
    output px2920 ;
    input \p_Pc_Add4(9)   ;
    output px2918 ;
    input \p_Pc_Add4(8)   ;
    output px2916 ;
    input \p_Pc_Add4(7)   ;
    output px2914 ;
    input \p_Pc_Add4(6)   ;
    output px2912 ;
    input \p_Pc_Add4(5)   ;
    output px2910 ;
    input \p_Pc_Add4(4)   ;
    output px2908 ;
    input \p_Pc_Add4(3)   ;
    output px2906 ;
    input \p_Pc_Add4(2)   ;
    output px2904 ;
    input [31:30]p_nbus_Addr_1_0 ;
    output px2902 ;
    input p_Ex_Z ;
    output px2900 ;
    input \p_Rt_1_0(2)   ;
    input \p_Rt_1_0(1)   ;
    input \p_Rt_1_0(0)   ;
    input \p_Id_Extimm(0)   ;
    output \p_Ex_Extimm(0)   ;
    input \p_Id_Extimm(1)   ;
    input \p_Id_Extimm(2)   ;
    input \p_Id_Extimm(3)   ;
    input \p_Id_Extimm(4)   ;
    input \p_Id_Extimm(13)   ;
    output \p_Ex_Extimm(13)   ;
    input \p_Id_Inst(26)   ;
    output \p_Ex_Op(0)   ;
    input \p_Id_Extimm(11)   ;
    input \p_Id_Extimm(12)   ;
    input \p_Id_Inst(28)   ;
    input \p_Id_Inst(29)   ;
    output [2:0]p_nbus_Ex_Rd ;
    output [2:0]p_nbus_Ex_Aluc ;
    input px3253 ;
    output [1:0]p_nbus_Ex_Fwd_A ;
    output px3255 ;
    input px3256 ;
    output [1:0]p_nbus_Ex_Fwd_B ;
    output px3258 ;
    output p_Ex_Wreg ;
    output p_Ex_Reg2reg ;
    output p_Ex_Wmem ;
    output p_Ex_Aluqb ;
    input [31:0]p_nbus_Id_Pc_Add4 ;
    output px3444 ;
    input p_EN_int ;
    input p_CLK_int ;
    input px2857 ;

    wire nx15296z4, nx15296z3, nx44340z2, nx45337z3, nx45337z2, \Ex_Extimm(1)  , 
         \Ex_Extimm(2)  , \Ex_Extimm(3)  , \Ex_Extimm(4)  , \Ex_Extimm(11)  , 
         \Ex_Extimm(12)  , \Ex_Op(2)  , \Ex_Op(3)  , nx19892z1, nx20889z1, 
         nx21886z1, nx45337z1, nx44340z1, nx43343z1, nx35354z1, nx10413z1, 
         nx24657z1, nx31806z1;
    wire [31:0]Ex_Pc;
    wire \Ex_Pc_0n1s1(31)  , nx36549z1, \Ex_Pc_0n1s1(30)  , nx36549z2, 
         \Ex_Pc_0n1s1(29)  , nx36549z3, \Ex_Pc_0n1s1(28)  , nx36549z4, 
         \Ex_Pc_0n1s1(27)  , nx36549z5, \Ex_Pc_0n1s1(26)  , nx36549z6, 
         \Ex_Pc_0n1s1(25)  , nx36549z7, \Ex_Pc_0n1s1(24)  , nx36549z8, 
         \Ex_Pc_0n1s1(23)  , nx36549z9, \Ex_Pc_0n1s1(22)  , nx36549z10, 
         \Ex_Pc_0n1s1(21)  , nx36549z11, \Ex_Pc_0n1s1(20)  , nx36549z12, 
         \Ex_Pc_0n1s1(19)  , nx36549z13, \Ex_Pc_0n1s1(18)  , nx36549z14, 
         \Ex_Pc_0n1s1(17)  , nx36549z15, \Ex_Pc_0n1s1(16)  , nx36549z16, 
         nx36549z40, \Ex_Pc_0n1s1(15)  , nx36549z17, nx36549z39, 
         \Ex_Pc_0n1s1(14)  , nx36549z18, nx36549z38, \Ex_Pc_0n1s1(13)  , 
         nx36549z19, \Ex_Pc_0n1s1(12)  , nx36549z20, \Ex_Pc_0n1s1(11)  , 
         nx36549z21, \Ex_Pc_0n1s1(10)  , nx36549z22, \Ex_Pc_0n1s1(9)  , 
         nx36549z23, nx36549z37, \Ex_Pc_0n1s1(8)  , nx36549z24, nx36549z36, 
         \Ex_Pc_0n1s1(7)  , nx36549z25, nx36549z35, \Ex_Pc_0n1s1(6)  , 
         nx36549z26, nx36549z34, \Ex_Pc_0n1s1(5)  , nx36549z27, nx36549z33, 
         \Ex_Pc_0n1s1(4)  , nx36549z28, nx36549z32, \Ex_Pc_0n1s1(3)  , 
         nx36549z29, nx36549z31, \Ex_Pc_0n1s1(2)  ;



    XORCY ix40575z19564 (.O (\Ex_Pc_0n1s1(2)  ), .CI (px2857), .LI (nx36549z31)
          ) ;
    XORCY ix41572z19564 (.O (\Ex_Pc_0n1s1(3)  ), .CI (nx36549z29), .LI (
          nx36549z32)) ;
    XORCY ix42569z19564 (.O (\Ex_Pc_0n1s1(4)  ), .CI (nx36549z28), .LI (
          nx36549z33)) ;
    XORCY ix43566z19564 (.O (\Ex_Pc_0n1s1(5)  ), .CI (nx36549z27), .LI (
          nx36549z34)) ;
    XORCY ix44563z19564 (.O (\Ex_Pc_0n1s1(6)  ), .CI (nx36549z26), .LI (
          nx36549z35)) ;
    XORCY ix45560z19564 (.O (\Ex_Pc_0n1s1(7)  ), .CI (nx36549z25), .LI (
          nx36549z36)) ;
    XORCY ix46557z19564 (.O (\Ex_Pc_0n1s1(8)  ), .CI (nx36549z24), .LI (
          nx36549z37)) ;
    XORCY ix47554z19564 (.O (\Ex_Pc_0n1s1(9)  ), .CI (nx36549z23), .LI (
          p_nbus_Id_Pc_Add4[7])) ;
    XORCY ix13614z19564 (.O (\Ex_Pc_0n1s1(10)  ), .CI (nx36549z22), .LI (
          p_nbus_Id_Pc_Add4[8])) ;
    XORCY ix14611z19564 (.O (\Ex_Pc_0n1s1(11)  ), .CI (nx36549z21), .LI (
          p_nbus_Id_Pc_Add4[9])) ;
    XORCY ix15608z19564 (.O (\Ex_Pc_0n1s1(12)  ), .CI (nx36549z20), .LI (
          p_nbus_Id_Pc_Add4[10])) ;
    XORCY ix16605z19564 (.O (\Ex_Pc_0n1s1(13)  ), .CI (nx36549z19), .LI (
          nx36549z38)) ;
    XORCY ix17602z19564 (.O (\Ex_Pc_0n1s1(14)  ), .CI (nx36549z18), .LI (
          nx36549z39)) ;
    XORCY ix18599z19564 (.O (\Ex_Pc_0n1s1(15)  ), .CI (nx36549z17), .LI (
          nx36549z40)) ;
    XORCY ix19596z19564 (.O (\Ex_Pc_0n1s1(16)  ), .CI (nx36549z16), .LI (
          p_nbus_Id_Pc_Add4[14])) ;
    XORCY ix20593z19564 (.O (\Ex_Pc_0n1s1(17)  ), .CI (nx36549z15), .LI (
          p_nbus_Id_Pc_Add4[15])) ;
    XORCY ix21590z19564 (.O (\Ex_Pc_0n1s1(18)  ), .CI (nx36549z14), .LI (
          p_nbus_Id_Pc_Add4[16])) ;
    XORCY ix22587z19564 (.O (\Ex_Pc_0n1s1(19)  ), .CI (nx36549z13), .LI (
          p_nbus_Id_Pc_Add4[17])) ;
    XORCY ix24583z19564 (.O (\Ex_Pc_0n1s1(20)  ), .CI (nx36549z12), .LI (
          p_nbus_Id_Pc_Add4[18])) ;
    XORCY ix25580z19564 (.O (\Ex_Pc_0n1s1(21)  ), .CI (nx36549z11), .LI (
          p_nbus_Id_Pc_Add4[19])) ;
    XORCY ix26577z19564 (.O (\Ex_Pc_0n1s1(22)  ), .CI (nx36549z10), .LI (
          p_nbus_Id_Pc_Add4[20])) ;
    XORCY ix27574z19564 (.O (\Ex_Pc_0n1s1(23)  ), .CI (nx36549z9), .LI (
          p_nbus_Id_Pc_Add4[21])) ;
    XORCY ix28571z19564 (.O (\Ex_Pc_0n1s1(24)  ), .CI (nx36549z8), .LI (
          p_nbus_Id_Pc_Add4[22])) ;
    XORCY ix29568z19564 (.O (\Ex_Pc_0n1s1(25)  ), .CI (nx36549z7), .LI (
          p_nbus_Id_Pc_Add4[23])) ;
    XORCY ix30565z19564 (.O (\Ex_Pc_0n1s1(26)  ), .CI (nx36549z6), .LI (
          p_nbus_Id_Pc_Add4[24])) ;
    XORCY ix31562z19564 (.O (\Ex_Pc_0n1s1(27)  ), .CI (nx36549z5), .LI (
          p_nbus_Id_Pc_Add4[25])) ;
    XORCY ix32559z19564 (.O (\Ex_Pc_0n1s1(28)  ), .CI (nx36549z4), .LI (
          p_nbus_Id_Pc_Add4[26])) ;
    XORCY ix33556z19564 (.O (\Ex_Pc_0n1s1(29)  ), .CI (nx36549z3), .LI (
          p_nbus_Id_Pc_Add4[27])) ;
    XORCY ix35552z19564 (.O (\Ex_Pc_0n1s1(30)  ), .CI (nx36549z2), .LI (
          p_nbus_Id_Pc_Add4[28])) ;
    XORCY ix36549z19564 (.O (\Ex_Pc_0n1s1(31)  ), .CI (nx36549z1), .LI (
          p_nbus_Id_Pc_Add4[29])) ;
    FDRE \reg_Ex_Pc(31)  (.Q (Ex_Pc[31]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(31)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(30)  (.Q (Ex_Pc[30]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(30)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(29)  (.Q (Ex_Pc[29]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(29)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(28)  (.Q (Ex_Pc[28]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(28)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(27)  (.Q (Ex_Pc[27]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(27)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(26)  (.Q (Ex_Pc[26]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(26)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(25)  (.Q (Ex_Pc[25]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(25)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(24)  (.Q (Ex_Pc[24]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(24)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(23)  (.Q (Ex_Pc[23]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(23)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(22)  (.Q (Ex_Pc[22]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(22)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(21)  (.Q (Ex_Pc[21]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(21)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(20)  (.Q (Ex_Pc[20]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(20)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(19)  (.Q (Ex_Pc[19]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(19)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(18)  (.Q (Ex_Pc[18]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(18)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(17)  (.Q (Ex_Pc[17]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(17)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(16)  (.Q (Ex_Pc[16]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(16)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(15)  (.Q (Ex_Pc[15]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(15)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(14)  (.Q (Ex_Pc[14]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(14)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(13)  (.Q (Ex_Pc[13]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(13)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(12)  (.Q (Ex_Pc[12]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(12)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(11)  (.Q (Ex_Pc[11]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(11)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(10)  (.Q (Ex_Pc[10]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(10)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(9)  (.Q (Ex_Pc[9]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(9)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(8)  (.Q (Ex_Pc[8]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(8)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(7)  (.Q (Ex_Pc[7]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(7)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(6)  (.Q (Ex_Pc[6]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(6)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(5)  (.Q (Ex_Pc[5]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(5)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(4)  (.Q (Ex_Pc[4]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(4)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(3)  (.Q (Ex_Pc[3]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(3)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(2)  (.Q (Ex_Pc[2]), .C (p_CLK_int), .CE (p_EN_int), .D (
         \Ex_Pc_0n1s1(2)  ), .R (px3444)) ;
    FDRE \reg_Ex_Pc(1)  (.Q (Ex_Pc[1]), .C (p_CLK_int), .CE (p_EN_int), .D (
         p_nbus_Id_Pc_Add4[30]), .R (px3444)) ;
    FDRE \reg_Ex_Pc(0)  (.Q (Ex_Pc[0]), .C (p_CLK_int), .CE (p_EN_int), .D (
         p_nbus_Id_Pc_Add4[31]), .R (px3444)) ;
    FDRE reg_Ex_Aluqb (.Q (p_Ex_Aluqb), .C (p_CLK_int), .CE (p_EN_int), .D (
         nx31806z1), .R (px3444)) ;
    FDRE reg_Ex_Wmem (.Q (p_Ex_Wmem), .C (p_CLK_int), .CE (p_EN_int), .D (
         nx24657z1), .R (px3444)) ;
    FDRE reg_Ex_Reg2reg (.Q (p_Ex_Reg2reg), .C (p_CLK_int), .CE (p_EN_int), .D (
         nx10413z1), .R (px3444)) ;
    FDRE reg_Ex_Wreg (.Q (p_Ex_Wreg), .C (p_CLK_int), .CE (p_EN_int), .D (
         nx35354z1), .R (px3444)) ;
    FDRE \reg_Ex_Fwd_B(1)  (.Q (p_nbus_Ex_Fwd_B[0]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3258), .R (px3444)) ;
    FDRE \reg_Ex_Fwd_B(0)  (.Q (p_nbus_Ex_Fwd_B[1]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3256), .R (px3444)) ;
    FDRE \reg_Ex_Fwd_A(1)  (.Q (p_nbus_Ex_Fwd_A[0]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3255), .R (px3444)) ;
    FDRE \reg_Ex_Fwd_A(0)  (.Q (p_nbus_Ex_Fwd_A[1]), .C (p_CLK_int), .CE (
         p_EN_int), .D (px3253), .R (px3444)) ;
    FDRE \reg_Ex_Aluc(2)  (.Q (p_nbus_Ex_Aluc[0]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (nx43343z1), .R (px3444)) ;
    FDRE \reg_Ex_Aluc(1)  (.Q (p_nbus_Ex_Aluc[1]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (nx44340z1), .R (px3444)) ;
    FDRE \reg_Ex_Aluc(0)  (.Q (p_nbus_Ex_Aluc[2]), .C (p_CLK_int), .CE (p_EN_int
         ), .D (nx45337z1), .R (px3444)) ;
    FDRE \reg_Ex_Rd(2)  (.Q (p_nbus_Ex_Rd[0]), .C (p_CLK_int), .CE (p_EN_int), .D (
         nx21886z1), .R (px3444)) ;
    FDRE \reg_Ex_Rd(1)  (.Q (p_nbus_Ex_Rd[1]), .C (p_CLK_int), .CE (p_EN_int), .D (
         nx20889z1), .R (px3444)) ;
    FDRE \reg_Ex_Rd(0)  (.Q (p_nbus_Ex_Rd[2]), .C (p_CLK_int), .CE (p_EN_int), .D (
         nx19892z1), .R (px3444)) ;
    FDRE \reg_Ex_Op(3)  (.Q (\Ex_Op(3)  ), .C (p_CLK_int), .CE (p_EN_int), .D (
         \p_Id_Inst(29)  ), .R (px3444)) ;
    FDRE \reg_Ex_Op(2)  (.Q (\Ex_Op(2)  ), .C (p_CLK_int), .CE (p_EN_int), .D (
         \p_Id_Inst(28)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(12)  (.Q (\Ex_Extimm(12)  ), .C (p_CLK_int), .CE (
         p_EN_int), .D (\p_Id_Extimm(12)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(11)  (.Q (\Ex_Extimm(11)  ), .C (p_CLK_int), .CE (
         p_EN_int), .D (\p_Id_Extimm(11)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(6)  (.Q (\p_Ex_Op(0)  ), .C (p_CLK_int), .CE (p_EN_int)
         , .D (\p_Id_Inst(26)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(5)  (.Q (\p_Ex_Extimm(13)  ), .C (p_CLK_int), .CE (
         p_EN_int), .D (\p_Id_Extimm(13)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(4)  (.Q (\Ex_Extimm(4)  ), .C (p_CLK_int), .CE (p_EN_int
         ), .D (\p_Id_Extimm(4)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(3)  (.Q (\Ex_Extimm(3)  ), .C (p_CLK_int), .CE (p_EN_int
         ), .D (\p_Id_Extimm(3)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(2)  (.Q (\Ex_Extimm(2)  ), .C (p_CLK_int), .CE (p_EN_int
         ), .D (\p_Id_Extimm(2)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(1)  (.Q (\Ex_Extimm(1)  ), .C (p_CLK_int), .CE (p_EN_int
         ), .D (\p_Id_Extimm(1)  ), .R (px3444)) ;
    FDRE \reg_Ex_Extimm(0)  (.Q (\p_Ex_Extimm(0)  ), .C (p_CLK_int), .CE (
         p_EN_int), .D (\p_Id_Extimm(0)  ), .R (px3444)) ;
    (* HLUTNM = "LUT62_3_2" *)
    LUT5 ix19892z45002 (.O (nx19892z1), .I0 (\p_Rt_1_0(0)  ), .I1 (
         \p_Id_Inst(29)  ), .I2 (\p_Id_Inst(28)  ), .I3 (\p_Id_Inst(26)  ), .I4 (
         \p_Id_Extimm(11)  )) ;
         defparam ix19892z45002.INIT = 32'hAAABAAA8;
    (* HLUTNM = "LUT62_3_3" *)
    LUT5 ix20889z45002 (.O (nx20889z1), .I0 (\p_Rt_1_0(1)  ), .I1 (
         \p_Id_Inst(29)  ), .I2 (\p_Id_Inst(28)  ), .I3 (\p_Id_Inst(26)  ), .I4 (
         \p_Id_Extimm(12)  )) ;
         defparam ix20889z45002.INIT = 32'hAAABAAA8;
    (* HLUTNM = "LUT62_3_4" *)
    LUT5 ix21886z45002 (.O (nx21886z1), .I0 (\p_Rt_1_0(2)  ), .I1 (
         \p_Id_Inst(29)  ), .I2 (\p_Id_Inst(28)  ), .I3 (\p_Id_Inst(26)  ), .I4 (
         \p_Id_Extimm(13)  )) ;
         defparam ix21886z45002.INIT = 32'hAAABAAA8;
    (* HLUTNM = "LUT62_3_2" *)
    LUT3 ix10413z1553 (.O (nx10413z1), .I0 (\p_Id_Inst(29)  ), .I1 (
         \p_Id_Inst(28)  ), .I2 (\p_Id_Inst(26)  )) ;
         defparam ix10413z1553.INIT = 8'hEF;
    (* HLUTNM = "LUT62_3_4" *)
    LUT3 ix31806z1511 (.O (nx31806z1), .I0 (\p_Id_Inst(29)  ), .I1 (
         \p_Id_Inst(28)  ), .I2 (\p_Id_Inst(26)  )) ;
         defparam ix31806z1511.INIT = 8'hC5;
    LUT2 ix36549z1359 (.O (nx36549z40), .I0 (p_nbus_Id_Pc_Add4[13]), .I1 (
         \p_Id_Extimm(13)  )) ;
         defparam ix36549z1359.INIT = 4'h6;
    LUT2 ix36549z1358 (.O (nx36549z39), .I0 (p_nbus_Id_Pc_Add4[12]), .I1 (
         \p_Id_Extimm(12)  )) ;
         defparam ix36549z1358.INIT = 4'h6;
    LUT2 ix36549z1357 (.O (nx36549z38), .I0 (p_nbus_Id_Pc_Add4[11]), .I1 (
         \p_Id_Extimm(11)  )) ;
         defparam ix36549z1357.INIT = 4'h6;
    LUT2 ix36549z1356 (.O (nx36549z37), .I0 (p_nbus_Id_Pc_Add4[6]), .I1 (
         \p_Id_Inst(26)  )) ;
         defparam ix36549z1356.INIT = 4'h6;
    LUT2 ix36549z1355 (.O (nx36549z36), .I0 (p_nbus_Id_Pc_Add4[5]), .I1 (
         \p_Id_Extimm(13)  )) ;
         defparam ix36549z1355.INIT = 4'h6;
    LUT2 ix36549z1354 (.O (nx36549z35), .I0 (p_nbus_Id_Pc_Add4[4]), .I1 (
         \p_Id_Extimm(4)  )) ;
         defparam ix36549z1354.INIT = 4'h6;
    LUT2 ix36549z1353 (.O (nx36549z34), .I0 (p_nbus_Id_Pc_Add4[3]), .I1 (
         \p_Id_Extimm(3)  )) ;
         defparam ix36549z1353.INIT = 4'h6;
    LUT2 ix36549z1352 (.O (nx36549z33), .I0 (p_nbus_Id_Pc_Add4[2]), .I1 (
         \p_Id_Extimm(2)  )) ;
         defparam ix36549z1352.INIT = 4'h6;
    LUT2 ix36549z1351 (.O (nx36549z32), .I0 (p_nbus_Id_Pc_Add4[1]), .I1 (
         \p_Id_Extimm(1)  )) ;
         defparam ix36549z1351.INIT = 4'h6;
    LUT2 ix36549z1350 (.O (nx36549z31), .I0 (p_nbus_Id_Pc_Add4[0]), .I1 (
         \p_Id_Extimm(0)  )) ;
         defparam ix36549z1350.INIT = 4'h6;
    LUT6 ix56509z45004 (.O (px2900), .I0 (p_nbus_Addr_1_0[30]), .I1 (Ex_Pc[0]), 
         .I2 (\Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)
         ) ;
         defparam ix56509z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix56507z45004 (.O (px2902), .I0 (p_nbus_Addr_1_0[31]), .I1 (Ex_Pc[1]), 
         .I2 (\Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)
         ) ;
         defparam ix56507z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix56505z45004 (.O (px2904), .I0 (\p_Pc_Add4(2)  ), .I1 (Ex_Pc[2]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix56505z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix56503z45004 (.O (px2906), .I0 (\p_Pc_Add4(3)  ), .I1 (Ex_Pc[3]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix56503z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix56501z45004 (.O (px2908), .I0 (\p_Pc_Add4(4)  ), .I1 (Ex_Pc[4]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix56501z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix55512z45004 (.O (px2910), .I0 (\p_Pc_Add4(5)  ), .I1 (Ex_Pc[5]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix55512z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix55510z45004 (.O (px2912), .I0 (\p_Pc_Add4(6)  ), .I1 (Ex_Pc[6]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix55510z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix55508z45004 (.O (px2914), .I0 (\p_Pc_Add4(7)  ), .I1 (Ex_Pc[7]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix55508z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix55506z45004 (.O (px2916), .I0 (\p_Pc_Add4(8)  ), .I1 (Ex_Pc[8]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix55506z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix55504z45004 (.O (px2918), .I0 (\p_Pc_Add4(9)  ), .I1 (Ex_Pc[9]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix55504z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix54515z45004 (.O (px2920), .I0 (\p_Pc_Add4(10)  ), .I1 (Ex_Pc[10]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix54515z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix54513z45004 (.O (px2922), .I0 (\p_Pc_Add4(11)  ), .I1 (Ex_Pc[11]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix54513z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix54511z45004 (.O (px2924), .I0 (\p_Pc_Add4(12)  ), .I1 (Ex_Pc[12]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix54511z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix54509z45004 (.O (px2926), .I0 (\p_Pc_Add4(13)  ), .I1 (Ex_Pc[13]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix54509z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix54507z45004 (.O (px2928), .I0 (\p_Pc_Add4(14)  ), .I1 (Ex_Pc[14]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix54507z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix53518z45004 (.O (px2930), .I0 (\p_Pc_Add4(15)  ), .I1 (Ex_Pc[15]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix53518z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix53516z45004 (.O (px2932), .I0 (\p_Pc_Add4(16)  ), .I1 (Ex_Pc[16]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix53516z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix53514z45004 (.O (px2934), .I0 (\p_Pc_Add4(17)  ), .I1 (Ex_Pc[17]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix53514z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix53512z45004 (.O (px2936), .I0 (\p_Pc_Add4(18)  ), .I1 (Ex_Pc[18]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix53512z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix53510z45004 (.O (px2938), .I0 (\p_Pc_Add4(19)  ), .I1 (Ex_Pc[19]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix53510z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix52521z45004 (.O (px2940), .I0 (\p_Pc_Add4(20)  ), .I1 (Ex_Pc[20]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix52521z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix52519z45004 (.O (px2942), .I0 (\p_Pc_Add4(21)  ), .I1 (Ex_Pc[21]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix52519z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix52517z45004 (.O (px2944), .I0 (\p_Pc_Add4(22)  ), .I1 (Ex_Pc[22]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix52517z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix52515z45004 (.O (px2946), .I0 (\p_Pc_Add4(23)  ), .I1 (Ex_Pc[23]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix52515z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix52513z45004 (.O (px2948), .I0 (\p_Pc_Add4(24)  ), .I1 (Ex_Pc[24]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix52513z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix51524z45004 (.O (px2950), .I0 (\p_Pc_Add4(25)  ), .I1 (Ex_Pc[25]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix51524z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix51522z45004 (.O (px2952), .I0 (\p_Pc_Add4(26)  ), .I1 (Ex_Pc[26]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix51522z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix51520z45004 (.O (px2954), .I0 (\p_Pc_Add4(27)  ), .I1 (Ex_Pc[27]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix51520z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix51518z45004 (.O (px2956), .I0 (\p_Pc_Add4(28)  ), .I1 (Ex_Pc[28]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix51518z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix51516z45004 (.O (px2958), .I0 (\p_Pc_Add4(29)  ), .I1 (Ex_Pc[29]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix51516z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix50527z45004 (.O (px2960), .I0 (\p_Pc_Add4(30)  ), .I1 (Ex_Pc[30]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix50527z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix50525z45004 (.O (px2962), .I0 (\p_Pc_Add4(31)  ), .I1 (Ex_Pc[31]), .I2 (
         \Ex_Op(3)  ), .I3 (\Ex_Op(2)  ), .I4 (\p_Ex_Op(0)  ), .I5 (p_Ex_Z)) ;
         defparam ix50525z45004.INIT = 64'hAAAAACAAAAAAAAAA;
    LUT6 ix47531z23278 (.O (px2995), .I0 (px3343), .I1 (\p_Ex_Extimm(13)  ), .I2 (
         p_nbus_Mem_Alu_R[30]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix47531z23278.INIT = 64'h55CC55CCF5CC55CC;
    LUT6 ix47530z542 (.O (px2996), .I0 (p_nbus_Ex_D2[26]), .I1 (\Ex_Extimm(12)  
         ), .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3347)) ;
         defparam ix47530z542.INIT = 64'hAC0C0CACFCFCFCFC;
    LUT6 ix47529z542 (.O (px2997), .I0 (p_nbus_Ex_D2[27]), .I1 (\Ex_Extimm(11)  
         ), .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3351)) ;
         defparam ix47529z542.INIT = 64'hAC0C0CACFCFCFCFC;
    LUT6 ix47528z14610 (.O (px2998), .I0 (px3462), .I1 (px3439), .I2 (
         \p_Ex_Op(0)  ), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix47528z14610.INIT = 64'h33F077F033F033F0;
    LUT6 ix47527z23278 (.O (px2999), .I0 (px3432), .I1 (\p_Ex_Extimm(13)  ), .I2 (
         p_nbus_Mem_Alu_R[31]), .I3 (p_Ex_Aluqb), .I4 (p_nbus_Ex_Fwd_B[0]), .I5 (
         p_nbus_Ex_Fwd_B[1])) ;
         defparam ix47527z23278.INIT = 64'h55CC55CCF5CC55CC;
    LUT6 ix32959z542 (.O (px3000), .I0 (p_nbus_Ex_D2[28]), .I1 (\Ex_Extimm(4)  )
         , .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3428)) ;
         defparam ix32959z542.INIT = 64'hAC0C0CACFCFCFCFC;
    LUT6 ix32960z542 (.O (px3001), .I0 (p_nbus_Ex_D2[29]), .I1 (\Ex_Extimm(3)  )
         , .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3424)) ;
         defparam ix32960z542.INIT = 64'hAC0C0CACFCFCFCFC;
    LUT6 ix32961z542 (.O (px3002), .I0 (p_nbus_Ex_D2[30]), .I1 (\Ex_Extimm(2)  )
         , .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3420)) ;
         defparam ix32961z542.INIT = 64'hAC0C0CACFCFCFCFC;
    LUT6 ix32962z542 (.O (px3003), .I0 (p_nbus_Ex_D2[31]), .I1 (\Ex_Extimm(1)  )
         , .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3367)) ;
         defparam ix32962z542.INIT = 64'hAC0C0CACFCFCFCFC;
    LUT6 ix54903z38187 (.O (px3206), .I0 (px3431), .I1 (px3430), .I2 (px3427), .I3 (
         px3426), .I4 (px3423), .I5 (px3422)) ;
         defparam ix54903z38187.INIT = 64'h9009000000009009;
    (* HLUTNM = "LUT62_3_1" *)
    LUT5 ix45337z22131 (.O (nx45337z1), .I0 (nx45337z2), .I1 (nx45337z3), .I2 (
         \p_Id_Extimm(3)  ), .I3 (\p_Id_Extimm(2)  ), .I4 (\p_Id_Extimm(1)  )) ;
         defparam ix45337z22131.INIT = 32'h55155151;
    (* HLUTNM = "LUT62_3_5" *)
    LUT4 ix44340z1508 (.O (nx44340z1), .I0 (nx44340z2), .I1 (\p_Id_Inst(29)  ), 
         .I2 (\p_Id_Inst(28)  ), .I3 (\p_Id_Inst(26)  )) ;
         defparam ix44340z1508.INIT = 16'h00C2;
    LUT5 ix44340z1827 (.O (nx44340z2), .I0 (\p_Id_Extimm(13)  ), .I1 (
         \p_Id_Extimm(4)  ), .I2 (\p_Id_Extimm(3)  ), .I3 (\p_Id_Extimm(2)  ), .I4 (
         \p_Id_Extimm(1)  )) ;
         defparam ix44340z1827.INIT = 32'h00000200;
    (* HLUTNM = "LUT62_3_1" *)
    LUT4 ix43343z3362 (.O (nx43343z1), .I0 (nx45337z3), .I1 (\p_Id_Extimm(3)  )
         , .I2 (\p_Id_Extimm(2)  ), .I3 (\p_Id_Extimm(1)  )) ;
         defparam ix43343z3362.INIT = 16'h0800;
    LUT6 ix45337z1572 (.O (nx45337z3), .I0 (\p_Id_Inst(29)  ), .I1 (
         \p_Id_Inst(28)  ), .I2 (\p_Id_Inst(26)  ), .I3 (\p_Id_Extimm(13)  ), .I4 (
         \p_Id_Extimm(4)  ), .I5 (\p_Id_Extimm(0)  )) ;
         defparam ix45337z1572.INIT = 64'h0000000000000100;
    LUT5 ix59887z1314 (.O (px3255), .I0 (nx15296z3), .I1 (p_nbus_Ex_Rd[0]), .I2 (
         p_nbus_Ex_Rd[1]), .I3 (p_nbus_Ex_Rd[2]), .I4 (p_Ex_Wreg)) ;
         defparam ix59887z1314.INIT = 32'hAAA80000;
    LUT5 ix17689z1314 (.O (px3258), .I0 (nx15296z4), .I1 (p_nbus_Ex_Rd[0]), .I2 (
         p_nbus_Ex_Rd[1]), .I3 (p_nbus_Ex_Rd[2]), .I4 (p_Ex_Wreg)) ;
         defparam ix17689z1314.INIT = 32'hAAA80000;
    (* HLUTNM = "LUT62_3_5" *)
    LUT3 ix35354z1533 (.O (nx35354z1), .I0 (\p_Id_Inst(29)  ), .I1 (
         \p_Id_Inst(28)  ), .I2 (\p_Id_Inst(26)  )) ;
         defparam ix35354z1533.INIT = 8'hDB;
    (* HLUTNM = "LUT62_3_3" *)
    LUT3 ix24657z1346 (.O (nx24657z1), .I0 (\p_Id_Inst(29)  ), .I1 (
         \p_Id_Inst(28)  ), .I2 (\p_Id_Inst(26)  )) ;
         defparam ix24657z1346.INIT = 8'h20;
    LUT3 ix45337z1373 (.O (nx45337z2), .I0 (\p_Id_Inst(29)  ), .I1 (
         \p_Id_Inst(28)  ), .I2 (\p_Id_Inst(26)  )) ;
         defparam ix45337z1373.INIT = 8'h3A;
    LUT6 ix4324z2085 (.O (px3346), .I0 (p_nbus_Ex_D2[26]), .I1 (\Ex_Extimm(12)  
         ), .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3347)) ;
         defparam ix4324z2085.INIT = 64'h53F3F35303030303;
    LUT6 ix5315z2085 (.O (px3350), .I0 (p_nbus_Ex_D2[27]), .I1 (\Ex_Extimm(11)  
         ), .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3351)) ;
         defparam ix5315z2085.INIT = 64'h53F3F35303030303;
    LUT6 ix6318z2085 (.O (px3366), .I0 (p_nbus_Ex_D2[31]), .I1 (\Ex_Extimm(1)  )
         , .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3367)) ;
         defparam ix6318z2085.INIT = 64'h53F3F35303030303;
    LUT4 ix6321z58130 (.O (px3369), .I0 (px3371), .I1 (px3370), .I2 (
         \p_Ex_Extimm(0)  ), .I3 (p_Ex_Aluqb)) ;
         defparam ix6321z58130.INIT = 16'hDDF0;
    LUT6 ix12305z2085 (.O (px3419), .I0 (p_nbus_Ex_D2[30]), .I1 (\Ex_Extimm(2)  
         ), .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3420)) ;
         defparam ix12305z2085.INIT = 64'h53F3F35303030303;
    LUT6 ix13296z2085 (.O (px3423), .I0 (p_nbus_Ex_D2[29]), .I1 (\Ex_Extimm(3)  
         ), .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3424)) ;
         defparam ix13296z2085.INIT = 64'h53F3F35303030303;
    LUT6 ix13300z2085 (.O (px3427), .I0 (p_nbus_Ex_D2[28]), .I1 (\Ex_Extimm(4)  
         ), .I2 (p_Ex_Aluqb), .I3 (p_nbus_Ex_Fwd_B[0]), .I4 (p_nbus_Ex_Fwd_B[1])
         , .I5 (px3428)) ;
         defparam ix13300z2085.INIT = 64'h53F3F35303030303;
    LUT4 ix21886z58899 (.O (px3444), .I0 (px3452), .I1 (px3450), .I2 (p_EN_int)
         , .I3 (p_CLR_N_int)) ;
         defparam ix21886z58899.INIT = 16'hE0F0;
    LUT4 ix15296z17778 (.O (px3449), .I0 (px3452), .I1 (px3450), .I2 (p_EN_int)
         , .I3 (p_CLR_N_int)) ;
         defparam ix15296z17778.INIT = 16'h4050;
    LUT4 ix21886z2340 (.O (px3450), .I0 (\Ex_Op(3)  ), .I1 (\Ex_Op(2)  ), .I2 (
         \p_Ex_Op(0)  ), .I3 (p_Ex_Z)) ;
         defparam ix21886z2340.INIT = 16'h0400;
    LUT6 ix15296z62467 (.O (px3452), .I0 (nx15296z3), .I1 (nx15296z4), .I2 (
         p_nbus_Ex_Rd[0]), .I3 (p_nbus_Ex_Rd[1]), .I4 (p_nbus_Ex_Rd[2]), .I5 (
         p_Ex_Reg2reg)) ;
         defparam ix15296z62467.INIT = 64'h00000000EEEEEEE0;
    LUT6 ix15296z1830 (.O (nx15296z4), .I0 (\p_Rt_1_0(2)  ), .I1 (\p_Rt_1_0(1)  
         ), .I2 (\p_Rt_1_0(0)  ), .I3 (p_nbus_Ex_Rd[0]), .I4 (p_nbus_Ex_Rd[1]), 
         .I5 (p_nbus_Ex_Rd[2])) ;
         defparam ix15296z1830.INIT = 64'h8040201008040201;
    LUT6 ix15296z1829 (.O (nx15296z3), .I0 (\p_Rs_1_0(2)  ), .I1 (\p_Rs_1_0(1)  
         ), .I2 (\p_Rs_1_0(0)  ), .I3 (p_nbus_Ex_Rd[0]), .I4 (p_nbus_Ex_Rd[1]), 
         .I5 (p_nbus_Ex_Rd[2])) ;
         defparam ix15296z1829.INIT = 64'h8040201008040201;
    MUXCY ix36549z63369 (.O (nx36549z29), .CI (px2857), .DI (
          p_nbus_Id_Pc_Add4[0]), .S (nx36549z31)) ;
    MUXCY ix36549z63368 (.O (nx36549z28), .CI (nx36549z29), .DI (
          p_nbus_Id_Pc_Add4[1]), .S (nx36549z32)) ;
    MUXCY ix36549z63367 (.O (nx36549z27), .CI (nx36549z28), .DI (
          p_nbus_Id_Pc_Add4[2]), .S (nx36549z33)) ;
    MUXCY ix36549z63366 (.O (nx36549z26), .CI (nx36549z27), .DI (
          p_nbus_Id_Pc_Add4[3]), .S (nx36549z34)) ;
    MUXCY ix36549z63365 (.O (nx36549z25), .CI (nx36549z26), .DI (
          p_nbus_Id_Pc_Add4[4]), .S (nx36549z35)) ;
    MUXCY ix36549z63364 (.O (nx36549z24), .CI (nx36549z25), .DI (
          p_nbus_Id_Pc_Add4[5]), .S (nx36549z36)) ;
    MUXCY ix36549z63363 (.O (nx36549z23), .CI (nx36549z24), .DI (
          p_nbus_Id_Pc_Add4[6]), .S (nx36549z37)) ;
    MUXCY ix36549z63362 (.O (nx36549z22), .CI (nx36549z23), .DI (
          p_nbus_Id_Pc_Add4[7]), .S (p_nbus_Id_Pc_Add4[7])) ;
    MUXCY ix36549z63361 (.O (nx36549z21), .CI (nx36549z22), .DI (
          p_nbus_Id_Pc_Add4[8]), .S (p_nbus_Id_Pc_Add4[8])) ;
    MUXCY ix36549z63360 (.O (nx36549z20), .CI (nx36549z21), .DI (
          p_nbus_Id_Pc_Add4[9]), .S (p_nbus_Id_Pc_Add4[9])) ;
    MUXCY ix36549z63359 (.O (nx36549z19), .CI (nx36549z20), .DI (
          p_nbus_Id_Pc_Add4[10]), .S (p_nbus_Id_Pc_Add4[10])) ;
    MUXCY ix36549z63358 (.O (nx36549z18), .CI (nx36549z19), .DI (
          p_nbus_Id_Pc_Add4[11]), .S (nx36549z38)) ;
    MUXCY ix36549z63357 (.O (nx36549z17), .CI (nx36549z18), .DI (
          p_nbus_Id_Pc_Add4[12]), .S (nx36549z39)) ;
    MUXCY ix36549z63356 (.O (nx36549z16), .CI (nx36549z17), .DI (
          p_nbus_Id_Pc_Add4[13]), .S (nx36549z40)) ;
    MUXCY ix36549z63355 (.O (nx36549z15), .CI (nx36549z16), .DI (
          p_nbus_Id_Pc_Add4[14]), .S (p_nbus_Id_Pc_Add4[14])) ;
    MUXCY ix36549z63354 (.O (nx36549z14), .CI (nx36549z15), .DI (
          p_nbus_Id_Pc_Add4[15]), .S (p_nbus_Id_Pc_Add4[15])) ;
    MUXCY ix36549z63353 (.O (nx36549z13), .CI (nx36549z14), .DI (
          p_nbus_Id_Pc_Add4[16]), .S (p_nbus_Id_Pc_Add4[16])) ;
    MUXCY ix36549z63352 (.O (nx36549z12), .CI (nx36549z13), .DI (
          p_nbus_Id_Pc_Add4[17]), .S (p_nbus_Id_Pc_Add4[17])) ;
    MUXCY ix36549z63351 (.O (nx36549z11), .CI (nx36549z12), .DI (
          p_nbus_Id_Pc_Add4[18]), .S (p_nbus_Id_Pc_Add4[18])) ;
    MUXCY ix36549z63350 (.O (nx36549z10), .CI (nx36549z11), .DI (
          p_nbus_Id_Pc_Add4[19]), .S (p_nbus_Id_Pc_Add4[19])) ;
    MUXCY ix36549z63349 (.O (nx36549z9), .CI (nx36549z10), .DI (
          p_nbus_Id_Pc_Add4[20]), .S (p_nbus_Id_Pc_Add4[20])) ;
    MUXCY ix36549z63348 (.O (nx36549z8), .CI (nx36549z9), .DI (
          p_nbus_Id_Pc_Add4[21]), .S (p_nbus_Id_Pc_Add4[21])) ;
    MUXCY ix36549z63347 (.O (nx36549z7), .CI (nx36549z8), .DI (
          p_nbus_Id_Pc_Add4[22]), .S (p_nbus_Id_Pc_Add4[22])) ;
    MUXCY ix36549z63346 (.O (nx36549z6), .CI (nx36549z7), .DI (
          p_nbus_Id_Pc_Add4[23]), .S (p_nbus_Id_Pc_Add4[23])) ;
    MUXCY ix36549z63345 (.O (nx36549z5), .CI (nx36549z6), .DI (
          p_nbus_Id_Pc_Add4[24]), .S (p_nbus_Id_Pc_Add4[24])) ;
    MUXCY ix36549z63344 (.O (nx36549z4), .CI (nx36549z5), .DI (
          p_nbus_Id_Pc_Add4[25]), .S (p_nbus_Id_Pc_Add4[25])) ;
    MUXCY ix36549z63343 (.O (nx36549z3), .CI (nx36549z4), .DI (
          p_nbus_Id_Pc_Add4[26]), .S (p_nbus_Id_Pc_Add4[26])) ;
    MUXCY ix36549z63342 (.O (nx36549z2), .CI (nx36549z3), .DI (
          p_nbus_Id_Pc_Add4[27]), .S (p_nbus_Id_Pc_Add4[27])) ;
    MUXCY ix36549z63341 (.O (nx36549z1), .CI (nx36549z2), .DI (
          p_nbus_Id_Pc_Add4[28]), .S (p_nbus_Id_Pc_Add4[28])) ;
endmodule


module REG_FILE_unfolded0_0 ( \p_Rs_1_0(0)  , \p_Rs_1_0(1)  , \p_Rs_1_0(2)  , 
                              \p_Rt_1_0(0)  , \p_Rt_1_0(1)  , \p_Rt_1_0(2)  , 
                              p_CLR_N_int, \p_Rd_1_0(0)  , \p_Rd_1_0(1)  , 
                              \p_Rd_1_0(2)  , p_rtlcs104, px3105, p_rtlcs103, 
                              px3104, p_rtlcs102, px3103, p_rtlcs101, px3102, 
                              p_rtlcs100, px3101, p_rtlcs99, px3100, p_rtlcs98, 
                              px3099, p_rtlcs97, px3098, p_rtlcs96, px3097, 
                              p_rtlcs95, px3096, p_rtlcs94, px3095, p_rtlcs93, 
                              px3094, p_rtlcs92, px3093, p_rtlcs91, px3092, 
                              p_rtlcs90, px3091, p_rtlcs89, px3090, p_rtlcs88, 
                              px3089, p_rtlcs87, px3088, p_rtlcs86, px3087, 
                              p_rtlcs85, px3086, p_rtlcs84, px3085, p_rtlcs83, 
                              px3084, p_rtlcs82, px3083, p_rtlcs81, px3082, 
                              p_rtlcs80, px3081, p_rtlcs79, px3080, p_rtlcs78, 
                              px3079, p_rtlcs77, px3078, p_rtlcs76, px3077, 
                              p_rtlcs75, px3076, p_rtlcs74, px3075, px3448, 
                              p_rtlcs73, px3074, p_rtlcs141, p_nbus_Wb_Alu_R, 
                              p_nbus_Wb_D, px3073, p_rtlcs140, px3072, 
                              p_rtlcs139, px3071, p_rtlcs138, px3070, p_rtlcs137, 
                              px3069, p_rtlcs136, px3068, p_rtlcs135, px3067, 
                              p_rtlcs134, px3066, p_rtlcs133, px3065, p_rtlcs132, 
                              px3064, p_rtlcs131, px3063, p_rtlcs130, px3062, 
                              p_rtlcs129, px3061, p_rtlcs128, px3060, p_rtlcs127, 
                              px3059, p_rtlcs126, px3058, p_rtlcs125, px3057, 
                              p_rtlcs124, px3056, p_rtlcs123, px3055, p_rtlcs122, 
                              px3054, p_rtlcs121, px3053, p_rtlcs120, px3052, 
                              p_rtlcs119, px3051, p_rtlcs118, px3050, p_rtlcs117, 
                              px3049, p_rtlcs116, px3048, p_rtlcs115, px3047, 
                              p_rtlcs114, px3046, p_rtlcs113, px3045, p_rtlcs112, 
                              px3044, p_rtlcs111, px3043, px3443, p_rtlcs110, 
                              p_Wb_Reg2reg, px3042, p_pc_not_clr_n, p_Wb_Wreg, 
                              p_CLK_int ) ;

    input \p_Rs_1_0(0)   ;
    input \p_Rs_1_0(1)   ;
    input \p_Rs_1_0(2)   ;
    input \p_Rt_1_0(0)   ;
    input \p_Rt_1_0(1)   ;
    input \p_Rt_1_0(2)   ;
    input p_CLR_N_int ;
    input \p_Rd_1_0(0)   ;
    input \p_Rd_1_0(1)   ;
    input \p_Rd_1_0(2)   ;
    input p_rtlcs104 ;
    output px3105 ;
    input p_rtlcs103 ;
    output px3104 ;
    input p_rtlcs102 ;
    output px3103 ;
    input p_rtlcs101 ;
    output px3102 ;
    input p_rtlcs100 ;
    output px3101 ;
    input p_rtlcs99 ;
    output px3100 ;
    input p_rtlcs98 ;
    output px3099 ;
    input p_rtlcs97 ;
    output px3098 ;
    input p_rtlcs96 ;
    output px3097 ;
    input p_rtlcs95 ;
    output px3096 ;
    input p_rtlcs94 ;
    output px3095 ;
    input p_rtlcs93 ;
    output px3094 ;
    input p_rtlcs92 ;
    output px3093 ;
    input p_rtlcs91 ;
    output px3092 ;
    input p_rtlcs90 ;
    output px3091 ;
    input p_rtlcs89 ;
    output px3090 ;
    input p_rtlcs88 ;
    output px3089 ;
    input p_rtlcs87 ;
    output px3088 ;
    input p_rtlcs86 ;
    output px3087 ;
    input p_rtlcs85 ;
    output px3086 ;
    input p_rtlcs84 ;
    output px3085 ;
    input p_rtlcs83 ;
    output px3084 ;
    input p_rtlcs82 ;
    output px3083 ;
    input p_rtlcs81 ;
    output px3082 ;
    input p_rtlcs80 ;
    output px3081 ;
    input p_rtlcs79 ;
    output px3080 ;
    input p_rtlcs78 ;
    output px3079 ;
    input p_rtlcs77 ;
    output px3078 ;
    input p_rtlcs76 ;
    output px3077 ;
    input p_rtlcs75 ;
    output px3076 ;
    input p_rtlcs74 ;
    output px3075 ;
    input px3448 ;
    input p_rtlcs73 ;
    output px3074 ;
    input p_rtlcs141 ;
    input [31:0]p_nbus_Wb_Alu_R ;
    input [31:0]p_nbus_Wb_D ;
    output px3073 ;
    input p_rtlcs140 ;
    output px3072 ;
    input p_rtlcs139 ;
    output px3071 ;
    input p_rtlcs138 ;
    output px3070 ;
    input p_rtlcs137 ;
    output px3069 ;
    input p_rtlcs136 ;
    output px3068 ;
    input p_rtlcs135 ;
    output px3067 ;
    input p_rtlcs134 ;
    output px3066 ;
    input p_rtlcs133 ;
    output px3065 ;
    input p_rtlcs132 ;
    output px3064 ;
    input p_rtlcs131 ;
    output px3063 ;
    input p_rtlcs130 ;
    output px3062 ;
    input p_rtlcs129 ;
    output px3061 ;
    input p_rtlcs128 ;
    output px3060 ;
    input p_rtlcs127 ;
    output px3059 ;
    input p_rtlcs126 ;
    output px3058 ;
    input p_rtlcs125 ;
    output px3057 ;
    input p_rtlcs124 ;
    output px3056 ;
    input p_rtlcs123 ;
    output px3055 ;
    input p_rtlcs122 ;
    output px3054 ;
    input p_rtlcs121 ;
    output px3053 ;
    input p_rtlcs120 ;
    output px3052 ;
    input p_rtlcs119 ;
    output px3051 ;
    input p_rtlcs118 ;
    output px3050 ;
    input p_rtlcs117 ;
    output px3049 ;
    input p_rtlcs116 ;
    output px3048 ;
    input p_rtlcs115 ;
    output px3047 ;
    input p_rtlcs114 ;
    output px3046 ;
    input p_rtlcs113 ;
    output px3045 ;
    input p_rtlcs112 ;
    output px3044 ;
    input p_rtlcs111 ;
    output px3043 ;
    input px3443 ;
    input p_rtlcs110 ;
    input p_Wb_Reg2reg ;
    output px3042 ;
    input p_pc_not_clr_n ;
    input p_Wb_Wreg ;
    input p_CLK_int ;

    wire nx43933z6, nx43933z5, nx39941z6, nx39941z5, nx43933z4, nx39941z4, 
         nx16240z1;
    wire [0:7]reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0;
    wire nx17237z1, nx18234z1, nx19231z1, nx20228z1, nx21225z1, nx22222z1, 
         nx23219z1, nx6, nx7, nx45, nx47, nx49, nx51, nx53, nx55, nx57;



    LUT6 ix36949z1314 (.O (px3042), .I0 (p_nbus_Wb_D[0]), .I1 (
         p_nbus_Wb_Alu_R[0]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs110), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36949z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix36950z1314 (.O (px3043), .I0 (p_nbus_Wb_D[1]), .I1 (
         p_nbus_Wb_Alu_R[1]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs111), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36950z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix36951z1314 (.O (px3044), .I0 (p_nbus_Wb_D[2]), .I1 (
         p_nbus_Wb_Alu_R[2]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs112), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36951z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix36952z1314 (.O (px3045), .I0 (p_nbus_Wb_D[3]), .I1 (
         p_nbus_Wb_Alu_R[3]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs113), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36952z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix36953z1314 (.O (px3046), .I0 (p_nbus_Wb_D[4]), .I1 (
         p_nbus_Wb_Alu_R[4]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs114), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36953z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix36954z1314 (.O (px3047), .I0 (p_nbus_Wb_D[5]), .I1 (
         p_nbus_Wb_Alu_R[5]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs115), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36954z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix36955z1314 (.O (px3048), .I0 (p_nbus_Wb_D[6]), .I1 (
         p_nbus_Wb_Alu_R[6]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs116), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36955z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix36956z1314 (.O (px3049), .I0 (p_nbus_Wb_D[7]), .I1 (
         p_nbus_Wb_Alu_R[7]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs117), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix36956z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37944z1314 (.O (px3050), .I0 (p_nbus_Wb_D[8]), .I1 (
         p_nbus_Wb_Alu_R[8]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs118), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix37944z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37945z1314 (.O (px3051), .I0 (p_nbus_Wb_D[9]), .I1 (
         p_nbus_Wb_Alu_R[9]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs119), .I4 (px3443)
         , .I5 (nx39941z4)) ;
         defparam ix37945z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37946z1314 (.O (px3052), .I0 (p_nbus_Wb_D[10]), .I1 (
         p_nbus_Wb_Alu_R[10]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs120), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37946z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37947z1314 (.O (px3053), .I0 (p_nbus_Wb_D[11]), .I1 (
         p_nbus_Wb_Alu_R[11]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs121), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37947z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37948z1314 (.O (px3054), .I0 (p_nbus_Wb_D[12]), .I1 (
         p_nbus_Wb_Alu_R[12]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs122), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37948z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37949z1314 (.O (px3055), .I0 (p_nbus_Wb_D[13]), .I1 (
         p_nbus_Wb_Alu_R[13]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs123), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37949z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37950z1314 (.O (px3056), .I0 (p_nbus_Wb_D[14]), .I1 (
         p_nbus_Wb_Alu_R[14]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs124), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37950z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37951z1314 (.O (px3057), .I0 (p_nbus_Wb_D[15]), .I1 (
         p_nbus_Wb_Alu_R[15]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs125), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37951z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37952z1314 (.O (px3058), .I0 (p_nbus_Wb_D[16]), .I1 (
         p_nbus_Wb_Alu_R[16]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs126), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37952z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix37953z1314 (.O (px3059), .I0 (p_nbus_Wb_D[17]), .I1 (
         p_nbus_Wb_Alu_R[17]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs127), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix37953z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38941z1314 (.O (px3060), .I0 (p_nbus_Wb_D[18]), .I1 (
         p_nbus_Wb_Alu_R[18]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs128), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38941z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38942z1314 (.O (px3061), .I0 (p_nbus_Wb_D[19]), .I1 (
         p_nbus_Wb_Alu_R[19]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs129), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38942z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38943z1314 (.O (px3062), .I0 (p_nbus_Wb_D[20]), .I1 (
         p_nbus_Wb_Alu_R[20]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs130), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38943z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38944z1314 (.O (px3063), .I0 (p_nbus_Wb_D[21]), .I1 (
         p_nbus_Wb_Alu_R[21]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs131), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38944z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38945z1314 (.O (px3064), .I0 (p_nbus_Wb_D[22]), .I1 (
         p_nbus_Wb_Alu_R[22]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs132), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38945z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38946z1314 (.O (px3065), .I0 (p_nbus_Wb_D[23]), .I1 (
         p_nbus_Wb_Alu_R[23]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs133), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38946z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38947z1314 (.O (px3066), .I0 (p_nbus_Wb_D[24]), .I1 (
         p_nbus_Wb_Alu_R[24]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs134), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38947z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38948z1314 (.O (px3067), .I0 (p_nbus_Wb_D[25]), .I1 (
         p_nbus_Wb_Alu_R[25]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs135), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38948z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38949z1314 (.O (px3068), .I0 (p_nbus_Wb_D[26]), .I1 (
         p_nbus_Wb_Alu_R[26]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs136), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38949z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix38950z1314 (.O (px3069), .I0 (p_nbus_Wb_D[27]), .I1 (
         p_nbus_Wb_Alu_R[27]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs137), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix38950z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39938z1314 (.O (px3070), .I0 (p_nbus_Wb_D[28]), .I1 (
         p_nbus_Wb_Alu_R[28]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs138), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix39938z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39939z1314 (.O (px3071), .I0 (p_nbus_Wb_D[29]), .I1 (
         p_nbus_Wb_Alu_R[29]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs139), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix39939z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39940z1314 (.O (px3072), .I0 (p_nbus_Wb_D[30]), .I1 (
         p_nbus_Wb_Alu_R[30]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs140), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix39940z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39941z1314 (.O (px3073), .I0 (p_nbus_Wb_D[31]), .I1 (
         p_nbus_Wb_Alu_R[31]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs141), .I4 (px3443
         ), .I5 (nx39941z4)) ;
         defparam ix39941z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39942z1314 (.O (px3074), .I0 (p_nbus_Wb_D[0]), .I1 (
         p_nbus_Wb_Alu_R[0]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs73), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix39942z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39943z1314 (.O (px3075), .I0 (p_nbus_Wb_D[1]), .I1 (
         p_nbus_Wb_Alu_R[1]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs74), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix39943z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39944z1314 (.O (px3076), .I0 (p_nbus_Wb_D[2]), .I1 (
         p_nbus_Wb_Alu_R[2]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs75), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix39944z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39945z1314 (.O (px3077), .I0 (p_nbus_Wb_D[3]), .I1 (
         p_nbus_Wb_Alu_R[3]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs76), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix39945z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39946z1314 (.O (px3078), .I0 (p_nbus_Wb_D[4]), .I1 (
         p_nbus_Wb_Alu_R[4]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs77), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix39946z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix39947z1314 (.O (px3079), .I0 (p_nbus_Wb_D[5]), .I1 (
         p_nbus_Wb_Alu_R[5]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs78), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix39947z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40935z1314 (.O (px3080), .I0 (p_nbus_Wb_D[6]), .I1 (
         p_nbus_Wb_Alu_R[6]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs79), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40935z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40936z1314 (.O (px3081), .I0 (p_nbus_Wb_D[7]), .I1 (
         p_nbus_Wb_Alu_R[7]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs80), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40936z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40937z1314 (.O (px3082), .I0 (p_nbus_Wb_D[8]), .I1 (
         p_nbus_Wb_Alu_R[8]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs81), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40937z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40938z1314 (.O (px3083), .I0 (p_nbus_Wb_D[9]), .I1 (
         p_nbus_Wb_Alu_R[9]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs82), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40938z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40939z1314 (.O (px3084), .I0 (p_nbus_Wb_D[10]), .I1 (
         p_nbus_Wb_Alu_R[10]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs83), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40939z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40940z1314 (.O (px3085), .I0 (p_nbus_Wb_D[11]), .I1 (
         p_nbus_Wb_Alu_R[11]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs84), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40940z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40941z1314 (.O (px3086), .I0 (p_nbus_Wb_D[12]), .I1 (
         p_nbus_Wb_Alu_R[12]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs85), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40941z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40942z1314 (.O (px3087), .I0 (p_nbus_Wb_D[13]), .I1 (
         p_nbus_Wb_Alu_R[13]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs86), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40942z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40943z1314 (.O (px3088), .I0 (p_nbus_Wb_D[14]), .I1 (
         p_nbus_Wb_Alu_R[14]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs87), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40943z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix40944z1314 (.O (px3089), .I0 (p_nbus_Wb_D[15]), .I1 (
         p_nbus_Wb_Alu_R[15]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs88), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix40944z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41932z1314 (.O (px3090), .I0 (p_nbus_Wb_D[16]), .I1 (
         p_nbus_Wb_Alu_R[16]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs89), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41932z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41933z1314 (.O (px3091), .I0 (p_nbus_Wb_D[17]), .I1 (
         p_nbus_Wb_Alu_R[17]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs90), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41933z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41934z1314 (.O (px3092), .I0 (p_nbus_Wb_D[18]), .I1 (
         p_nbus_Wb_Alu_R[18]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs91), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41934z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41935z1314 (.O (px3093), .I0 (p_nbus_Wb_D[19]), .I1 (
         p_nbus_Wb_Alu_R[19]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs92), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41935z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41936z1314 (.O (px3094), .I0 (p_nbus_Wb_D[20]), .I1 (
         p_nbus_Wb_Alu_R[20]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs93), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41936z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41937z1314 (.O (px3095), .I0 (p_nbus_Wb_D[21]), .I1 (
         p_nbus_Wb_Alu_R[21]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs94), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41937z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41938z1314 (.O (px3096), .I0 (p_nbus_Wb_D[22]), .I1 (
         p_nbus_Wb_Alu_R[22]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs95), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41938z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41939z1314 (.O (px3097), .I0 (p_nbus_Wb_D[23]), .I1 (
         p_nbus_Wb_Alu_R[23]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs96), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41939z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41940z1314 (.O (px3098), .I0 (p_nbus_Wb_D[24]), .I1 (
         p_nbus_Wb_Alu_R[24]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs97), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41940z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix41941z1314 (.O (px3099), .I0 (p_nbus_Wb_D[25]), .I1 (
         p_nbus_Wb_Alu_R[25]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs98), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix41941z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix43928z1314 (.O (px3100), .I0 (p_nbus_Wb_D[26]), .I1 (
         p_nbus_Wb_Alu_R[26]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs99), .I4 (px3448)
         , .I5 (nx43933z4)) ;
         defparam ix43928z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix43929z1314 (.O (px3101), .I0 (p_nbus_Wb_D[27]), .I1 (
         p_nbus_Wb_Alu_R[27]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs100), .I4 (px3448
         ), .I5 (nx43933z4)) ;
         defparam ix43929z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix43930z1314 (.O (px3102), .I0 (p_nbus_Wb_D[28]), .I1 (
         p_nbus_Wb_Alu_R[28]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs101), .I4 (px3448
         ), .I5 (nx43933z4)) ;
         defparam ix43930z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix43931z1314 (.O (px3103), .I0 (p_nbus_Wb_D[29]), .I1 (
         p_nbus_Wb_Alu_R[29]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs102), .I4 (px3448
         ), .I5 (nx43933z4)) ;
         defparam ix43931z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix43932z1314 (.O (px3104), .I0 (p_nbus_Wb_D[30]), .I1 (
         p_nbus_Wb_Alu_R[30]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs103), .I4 (px3448
         ), .I5 (nx43933z4)) ;
         defparam ix43932z1314.INIT = 64'hFFCAFF00CACA0000;
    LUT6 ix43933z1314 (.O (px3105), .I0 (p_nbus_Wb_D[31]), .I1 (
         p_nbus_Wb_Alu_R[31]), .I2 (p_Wb_Reg2reg), .I3 (p_rtlcs104), .I4 (px3448
         ), .I5 (nx43933z4)) ;
         defparam ix43933z1314.INIT = 64'hFFCAFF00CACA0000;
    (* HLUTNM = "LUT62_2_1" *)
    LUT5 ix16240z1314 (.O (nx16240z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix16240z1314.INIT = 32'h01000000;
    (* HLUTNM = "LUT62_2_1" *)
    LUT5 ix17237z1314 (.O (nx17237z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix17237z1314.INIT = 32'h10000000;
    (* HLUTNM = "LUT62_2_2" *)
    LUT5 ix18234z1314 (.O (nx18234z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix18234z1314.INIT = 32'h04000000;
    (* HLUTNM = "LUT62_2_2" *)
    LUT5 ix19231z1314 (.O (nx19231z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix19231z1314.INIT = 32'h40000000;
    (* HLUTNM = "LUT62_2_3" *)
    LUT5 ix20228z1314 (.O (nx20228z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix20228z1314.INIT = 32'h02000000;
    (* HLUTNM = "LUT62_2_3" *)
    LUT5 ix21225z1314 (.O (nx21225z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix21225z1314.INIT = 32'h20000000;
    (* HLUTNM = "LUT62_2_4" *)
    LUT5 ix22222z1314 (.O (nx22222z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix22222z1314.INIT = 32'h08000000;
    (* HLUTNM = "LUT62_2_4" *)
    LUT5 ix23219z1314 (.O (nx23219z1), .I0 (\p_Rd_1_0(2)  ), .I1 (\p_Rd_1_0(1)  
         ), .I2 (\p_Rd_1_0(0)  ), .I3 (p_Wb_Wreg), .I4 (p_CLR_N_int)) ;
         defparam ix23219z1314.INIT = 32'h80000000;
    LUT4 ix39941z18803 (.O (nx39941z4), .I0 (px3443), .I1 (nx39941z5), .I2 (
         nx39941z6), .I3 (\p_Rt_1_0(2)  )) ;
         defparam ix39941z18803.INIT = 16'h4450;
    LUT6 ix39941z45332 (.O (nx39941z6), .I0 (\p_Rt_1_0(1)  ), .I1 (\p_Rt_1_0(0)  
         ), .I2 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[0])
         , .I3 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[1])
         , .I4 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[2])
         , .I5 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[3])
         ) ;
         defparam ix39941z45332.INIT = 64'h0145236789CDABEF;
    LUT6 ix39941z45331 (.O (nx39941z5), .I0 (\p_Rt_1_0(1)  ), .I1 (\p_Rt_1_0(0)  
         ), .I2 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[4])
         , .I3 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[5])
         , .I4 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[6])
         , .I5 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[7])
         ) ;
         defparam ix39941z45331.INIT = 64'h0145236789CDABEF;
    LUT4 ix43933z18803 (.O (nx43933z4), .I0 (px3448), .I1 (nx43933z5), .I2 (
         nx43933z6), .I3 (\p_Rs_1_0(2)  )) ;
         defparam ix43933z18803.INIT = 16'h4450;
    LUT6 ix43933z45332 (.O (nx43933z6), .I0 (\p_Rs_1_0(1)  ), .I1 (\p_Rs_1_0(0)  
         ), .I2 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[0])
         , .I3 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[1])
         , .I4 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[2])
         , .I5 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[3])
         ) ;
         defparam ix43933z45332.INIT = 64'h0145236789CDABEF;
    LUT6 ix43933z45331 (.O (nx43933z5), .I0 (\p_Rs_1_0(1)  ), .I1 (\p_Rs_1_0(0)  
         ), .I2 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[4])
         , .I3 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[5])
         , .I4 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[6])
         , .I5 (reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[7])
         ) ;
         defparam ix43933z45331.INIT = 64'h0145236789CDABEF;
    VCC \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(7)_I21_FD_PWR  (
        .P (nx6)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(7)_I21_FD_LUT 
          (.O (nx7), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[7]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[7]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(7)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(7)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[7]), .C (
         p_CLK_int), .CE (nx6), .D (nx7), .R (nx23219z1)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(6)_I21_FD_LUT 
          (.O (nx45), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[6]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[6]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(6)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(6)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[6]), .C (
         p_CLK_int), .CE (nx6), .D (nx45), .R (nx22222z1)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(5)_I21_FD_LUT 
          (.O (nx47), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[5]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[5]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(5)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(5)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[5]), .C (
         p_CLK_int), .CE (nx6), .D (nx47), .R (nx21225z1)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(4)_I21_FD_LUT 
          (.O (nx49), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[4]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[4]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(4)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(4)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[4]), .C (
         p_CLK_int), .CE (nx6), .D (nx49), .R (nx20228z1)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(3)_I21_FD_LUT 
          (.O (nx51), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[3]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[3]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(3)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(3)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[3]), .C (
         p_CLK_int), .CE (nx6), .D (nx51), .R (nx19231z1)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(2)_I21_FD_LUT 
          (.O (nx53), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[2]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[2]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(2)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(2)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[2]), .C (
         p_CLK_int), .CE (nx6), .D (nx53), .R (nx18234z1)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(1)_I21_FD_LUT 
          (.O (nx55), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[1]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[1]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(1)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(1)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[1]), .C (
         p_CLK_int), .CE (nx6), .D (nx55), .R (nx17237z1)) ;
    LUT4 \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(0)_I21_FD_LUT 
          (.O (nx57), .I0 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[0]), .I1 (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[0]), .I2 (
         p_Wb_Wreg), .I3 (p_pc_not_clr_n)) ;
         defparam \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(0)_I21_FD_LUT .INIT = 16'hFFCA;
    FDRE \reg_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0(0)  (.Q (
         reg_file_MSR__REG_FILE_register_2_rtlc_sync_msr_n0_rtlcGen0[0]), .C (
         p_CLK_int), .CE (nx6), .D (nx57), .R (nx16240z1)) ;
endmodule


module INST_MEM_0 ( p_nbus_Addr_1_0, \p_Instruction(0)  , \p_Instruction(1)  , 
                    \p_Instruction(2)  , \p_Instruction(3)  , \p_Instruction(4)  , 
                    \p_Instruction(13)  , \p_Instruction(31)  , 
                    \p_Instruction(11)  , \p_Instruction(12)  , 
                    \p_Instruction(16)  , \p_Instruction(17)  , 
                    \p_Instruction(18)  , \p_Instruction(21)  , 
                    \p_Instruction(22)  , \p_Instruction(23)  , 
                    \p_Instruction(28)  , \p_Instruction(29)   ) ;

    input [31:0]p_nbus_Addr_1_0 ;
    output \p_Instruction(0)   ;
    output \p_Instruction(1)   ;
    output \p_Instruction(2)   ;
    output \p_Instruction(3)   ;
    output \p_Instruction(4)   ;
    output \p_Instruction(13)   ;
    output \p_Instruction(31)   ;
    output \p_Instruction(11)   ;
    output \p_Instruction(12)   ;
    output \p_Instruction(16)   ;
    output \p_Instruction(17)   ;
    output \p_Instruction(18)   ;
    output \p_Instruction(21)   ;
    output \p_Instruction(22)   ;
    output \p_Instruction(23)   ;
    output \p_Instruction(28)   ;
    output \p_Instruction(29)   ;

    wire nx33819z8, nx33819z7, nx33819z6, nx33819z5, nx33819z4, nx33819z10, 
         nx33819z9, nx33819z3, nx33819z1, nx34816z1, nx35813z1, nx36810z1, 
         nx37807z1, nx38804z1, nx39801z1, nx14511z1, nx13514z1, nx9526z1, 
         nx8529z1, nx7532z1, nx3542z1, nx2545z1, nx1548z1, nx62099z1, nx33819z2, 
         nx61102z1, nx3, nx4;



    (* HLUTNM = "LUT62_1_3" *)
    LUT5 ix35813z45021 (.O (nx35813z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix35813z45021.INIT = 32'hABEBAABB;
    (* HLUTNM = "LUT62_1_7" *)
    LUT4 ix36810z18050 (.O (nx36810z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix36810z18050.INIT = 16'h4160;
    (* HLUTNM = "LUT62_1_3" *)
    LUT5 ix37807z61388 (.O (nx37807z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix37807z61388.INIT = 32'hAAAAEAAA;
    (* HLUTNM = "LUT62_1_4" *)
    LUT5 ix39801z61388 (.O (nx39801z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix39801z61388.INIT = 32'hAAEAEAAA;
    (* HLUTNM = "LUT62_1_6" *)
    LUT4 ix14511z10542 (.O (nx14511z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix14511z10542.INIT = 16'h240C;
    (* HLUTNM = "LUT62_1_9" *)
    LUT4 ix9526z12402 (.O (nx9526z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix9526z12402.INIT = 16'h2B50;
    (* HLUTNM = "LUT62_1_5" *)
    LUT5 ix8529z1293 (.O (nx8529z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix8529z1293.INIT = 32'hEBEBFFEB;
    (* HLUTNM = "LUT62_1_9" *)
    LUT4 ix7532z29558 (.O (nx7532z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix7532z29558.INIT = 16'h6E54;
    (* HLUTNM = "LUT62_1_7" *)
    LUT4 ix3542z24974 (.O (nx3542z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix3542z24974.INIT = 16'h5C6C;
    (* HLUTNM = "LUT62_1_6" *)
    LUT4 ix2545z23886 (.O (nx2545z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix2545z23886.INIT = 16'h582C;
    (* HLUTNM = "LUT62_1_1" *)
    LUT5 ix33819z1575 (.O (nx33819z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix33819z1575.INIT = 32'h41000105;
    (* HLUTNM = "LUT62_1_2" *)
    LUT5 ix34816z6754 (.O (nx34816z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix34816z6754.INIT = 32'h10001540;
    (* HLUTNM = "LUT62_1_4" *)
    LUT5 ix38804z2418 (.O (nx38804z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix38804z2418.INIT = 32'h15100450;
    (* HLUTNM = "LUT62_1_5" *)
    LUT4 ix13514z9514 (.O (nx13514z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix13514z9514.INIT = 16'h2008;
    (* HLUTNM = "LUT62_1_1" *)
    LUT5 ix1548z6502 (.O (nx1548z1), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix1548z6502.INIT = 32'h05101444;
    (* HLUTNM = "LUT62_1_8" *)
    LUT4 ix62099z1380 (.O (nx62099z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix62099z1380.INIT = 16'h0042;
    LUT6 ix33819z1443 (.O (nx33819z2), .I0 (nx33819z3), .I1 (nx33819z9), .I2 (
         nx33819z10), .I3 (p_nbus_Addr_1_0[5]), .I4 (p_nbus_Addr_1_0[6]), .I5 (
         p_nbus_Addr_1_0[7])) ;
         defparam ix33819z1443.INIT = 64'h0000000000000080;
    LUT4 ix33819z1324 (.O (nx33819z10), .I0 (p_nbus_Addr_1_0[8]), .I1 (
         p_nbus_Addr_1_0[9]), .I2 (p_nbus_Addr_1_0[10]), .I3 (
         p_nbus_Addr_1_0[11])) ;
         defparam ix33819z1324.INIT = 16'h0001;
    LUT4 ix33819z1323 (.O (nx33819z9), .I0 (p_nbus_Addr_1_0[12]), .I1 (
         p_nbus_Addr_1_0[13]), .I2 (p_nbus_Addr_1_0[14]), .I3 (
         p_nbus_Addr_1_0[15])) ;
         defparam ix33819z1323.INIT = 16'h0001;
    LUT5 ix33819z34084 (.O (nx33819z3), .I0 (nx33819z4), .I1 (nx33819z5), .I2 (
         nx33819z6), .I3 (nx33819z7), .I4 (nx33819z8)) ;
         defparam ix33819z34084.INIT = 32'h00008000;
    (* HLUTNM = "LUT62_1_2" *)
    LUT5 ix33819z45009 (.O (nx33819z8), .I0 (p_nbus_Addr_1_0[0]), .I1 (
         p_nbus_Addr_1_0[1]), .I2 (p_nbus_Addr_1_0[2]), .I3 (p_nbus_Addr_1_0[3])
         , .I4 (p_nbus_Addr_1_0[4])) ;
         defparam ix33819z45009.INIT = 32'hAAAAAAA8;
    LUT4 ix33819z1321 (.O (nx33819z7), .I0 (p_nbus_Addr_1_0[16]), .I1 (
         p_nbus_Addr_1_0[17]), .I2 (p_nbus_Addr_1_0[18]), .I3 (
         p_nbus_Addr_1_0[19])) ;
         defparam ix33819z1321.INIT = 16'h0001;
    LUT4 ix33819z1320 (.O (nx33819z6), .I0 (p_nbus_Addr_1_0[20]), .I1 (
         p_nbus_Addr_1_0[21]), .I2 (p_nbus_Addr_1_0[22]), .I3 (
         p_nbus_Addr_1_0[23])) ;
         defparam ix33819z1320.INIT = 16'h0001;
    LUT4 ix33819z1319 (.O (nx33819z5), .I0 (p_nbus_Addr_1_0[24]), .I1 (
         p_nbus_Addr_1_0[25]), .I2 (p_nbus_Addr_1_0[26]), .I3 (
         p_nbus_Addr_1_0[27])) ;
         defparam ix33819z1319.INIT = 16'h0001;
    LUT4 ix33819z1318 (.O (nx33819z4), .I0 (p_nbus_Addr_1_0[28]), .I1 (
         p_nbus_Addr_1_0[29]), .I2 (p_nbus_Addr_1_0[30]), .I3 (
         p_nbus_Addr_1_0[31])) ;
         defparam ix33819z1318.INIT = 16'h0001;
    (* HLUTNM = "LUT62_1_8" *)
    LUT4 ix61102z36915 (.O (nx61102z1), .I0 (p_nbus_Addr_1_0[1]), .I1 (
         p_nbus_Addr_1_0[2]), .I2 (p_nbus_Addr_1_0[3]), .I3 (p_nbus_Addr_1_0[4])
         ) ;
         defparam ix61102z36915.INIT = 16'h8B11;
    VCC \lat_instruction(29)_I14_LD_PWR  (.P (nx3)) ;
    GND \lat_instruction(29)_I14_LD_GND  (.G (nx4)) ;
    LDCE \lat_instruction(29)  (.Q (\p_Instruction(29)  ), .CLR (nx4), .D (
         nx61102z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(28)  (.Q (\p_Instruction(28)  ), .CLR (nx4), .D (
         nx62099z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(23)  (.Q (\p_Instruction(23)  ), .CLR (nx4), .D (
         nx1548z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(22)  (.Q (\p_Instruction(22)  ), .CLR (nx4), .D (
         nx2545z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(21)  (.Q (\p_Instruction(21)  ), .CLR (nx4), .D (
         nx3542z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(18)  (.Q (\p_Instruction(18)  ), .CLR (nx4), .D (
         nx7532z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(17)  (.Q (\p_Instruction(17)  ), .CLR (nx4), .D (
         nx8529z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(16)  (.Q (\p_Instruction(16)  ), .CLR (nx4), .D (
         nx9526z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(12)  (.Q (\p_Instruction(12)  ), .CLR (nx4), .D (
         nx13514z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(11)  (.Q (\p_Instruction(11)  ), .CLR (nx4), .D (
         nx14511z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(6)  (.Q (\p_Instruction(31)  ), .CLR (nx4), .D (
         nx39801z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(5)  (.Q (\p_Instruction(13)  ), .CLR (nx4), .D (
         nx38804z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(4)  (.Q (\p_Instruction(4)  ), .CLR (nx4), .D (
         nx37807z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(3)  (.Q (\p_Instruction(3)  ), .CLR (nx4), .D (
         nx36810z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(2)  (.Q (\p_Instruction(2)  ), .CLR (nx4), .D (
         nx35813z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(1)  (.Q (\p_Instruction(1)  ), .CLR (nx4), .D (
         nx34816z1), .G (nx33819z2), .GE (nx3)) ;
    LDCE \lat_instruction(0)  (.Q (\p_Instruction(0)  ), .CLR (nx4), .D (
         nx33819z1), .G (nx33819z2), .GE (nx3)) ;
endmodule


module MUX4X32_0 ( px2900, p_nbus_Next_Addr, px2902, px2904, px2906, px2908, 
                   px2910, px2912, px2914, px2916, px2918, px2920, px2922, 
                   px2924, px2926, px2928, px2930, px2932, px2934, px2936, 
                   px2938, px2940, px2942, px2944, px2946, px2948, px2950, 
                   px2952, px2954, px2956, px2958, px2960, px2855, px2962 ) ;

    input px2900 ;
    output [31:0]p_nbus_Next_Addr ;
    input px2902 ;
    input px2904 ;
    input px2906 ;
    input px2908 ;
    input px2910 ;
    input px2912 ;
    input px2914 ;
    input px2916 ;
    input px2918 ;
    input px2920 ;
    input px2922 ;
    input px2924 ;
    input px2926 ;
    input px2928 ;
    input px2930 ;
    input px2932 ;
    input px2934 ;
    input px2936 ;
    input px2938 ;
    input px2940 ;
    input px2942 ;
    input px2944 ;
    input px2946 ;
    input px2948 ;
    input px2950 ;
    input px2952 ;
    input px2954 ;
    input px2956 ;
    input px2958 ;
    input px2960 ;
    input px2855 ;
    input px2962 ;

    wire nx3, nx4;



    VCC \lat_Out_addr(31)_I14_LD_PWR  (.P (nx3)) ;
    GND \lat_Out_addr(31)_I14_LD_GND  (.G (nx4)) ;
    LDCE \lat_Out_addr(31)  (.Q (p_nbus_Next_Addr[0]), .CLR (nx4), .D (px2962), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(30)  (.Q (p_nbus_Next_Addr[1]), .CLR (nx4), .D (px2960), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(29)  (.Q (p_nbus_Next_Addr[2]), .CLR (nx4), .D (px2958), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(28)  (.Q (p_nbus_Next_Addr[3]), .CLR (nx4), .D (px2956), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(27)  (.Q (p_nbus_Next_Addr[4]), .CLR (nx4), .D (px2954), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(26)  (.Q (p_nbus_Next_Addr[5]), .CLR (nx4), .D (px2952), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(25)  (.Q (p_nbus_Next_Addr[6]), .CLR (nx4), .D (px2950), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(24)  (.Q (p_nbus_Next_Addr[7]), .CLR (nx4), .D (px2948), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(23)  (.Q (p_nbus_Next_Addr[8]), .CLR (nx4), .D (px2946), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(22)  (.Q (p_nbus_Next_Addr[9]), .CLR (nx4), .D (px2944), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(21)  (.Q (p_nbus_Next_Addr[10]), .CLR (nx4), .D (px2942)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(20)  (.Q (p_nbus_Next_Addr[11]), .CLR (nx4), .D (px2940)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(19)  (.Q (p_nbus_Next_Addr[12]), .CLR (nx4), .D (px2938)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(18)  (.Q (p_nbus_Next_Addr[13]), .CLR (nx4), .D (px2936)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(17)  (.Q (p_nbus_Next_Addr[14]), .CLR (nx4), .D (px2934)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(16)  (.Q (p_nbus_Next_Addr[15]), .CLR (nx4), .D (px2932)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(15)  (.Q (p_nbus_Next_Addr[16]), .CLR (nx4), .D (px2930)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(14)  (.Q (p_nbus_Next_Addr[17]), .CLR (nx4), .D (px2928)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(13)  (.Q (p_nbus_Next_Addr[18]), .CLR (nx4), .D (px2926)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(12)  (.Q (p_nbus_Next_Addr[19]), .CLR (nx4), .D (px2924)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(11)  (.Q (p_nbus_Next_Addr[20]), .CLR (nx4), .D (px2922)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(10)  (.Q (p_nbus_Next_Addr[21]), .CLR (nx4), .D (px2920)
         , .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(9)  (.Q (p_nbus_Next_Addr[22]), .CLR (nx4), .D (px2918), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(8)  (.Q (p_nbus_Next_Addr[23]), .CLR (nx4), .D (px2916), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(7)  (.Q (p_nbus_Next_Addr[24]), .CLR (nx4), .D (px2914), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(6)  (.Q (p_nbus_Next_Addr[25]), .CLR (nx4), .D (px2912), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(5)  (.Q (p_nbus_Next_Addr[26]), .CLR (nx4), .D (px2910), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(4)  (.Q (p_nbus_Next_Addr[27]), .CLR (nx4), .D (px2908), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(3)  (.Q (p_nbus_Next_Addr[28]), .CLR (nx4), .D (px2906), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(2)  (.Q (p_nbus_Next_Addr[29]), .CLR (nx4), .D (px2904), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(1)  (.Q (p_nbus_Next_Addr[30]), .CLR (nx4), .D (px2902), 
         .G (px2855), .GE (nx3)) ;
    LDCE \lat_Out_addr(0)  (.Q (p_nbus_Next_Addr[31]), .CLR (nx4), .D (px2900), 
         .G (px2855), .GE (nx3)) ;
endmodule


module inc_30_0 ( cin, a, d, cout ) ;

    input cin ;
    input [29:0]a ;
    output [29:0]d ;
    output cout ;

    wire nx8473z2, nx8473z1, nx8473z3, nx8474z1, nx8474z2, nx8475z1, nx8475z2, 
         nx8476z1, nx8476z2, nx8477z1, nx8477z2, nx8478z1, nx8478z2, nx8479z1, 
         nx8479z2, nx8480z1, nx8480z2, nx8481z1, nx8481z2, nx8482z1, nx8482z2, 
         nx60018z1, nx60018z2, nx60019z1, nx60019z2, nx60020z1, nx60020z2, 
         nx60021z1, nx60021z2, nx60022z1, nx60022z2, nx60023z1, nx60023z2, 
         nx60024z1, nx60024z2, nx60025z1, nx60025z2, nx60026z1, nx60026z2, 
         nx60027z1, nx60027z2, nx61015z1, nx61015z2, nx61016z1, nx61016z2, 
         nx61017z1, nx61017z2, nx61018z1, nx61018z2, nx61019z1, nx61019z2, 
         nx61020z1, nx61020z2, nx61021z1, nx61021z2, nx61022z1, nx61022z2, 
         nx61023z1, nx61023z2, nx19589z1;



    GND ps_gnd (.G (nx8473z2)) ;
    VCC ps_vcc (.P (nx8473z1)) ;
    XORCY xorcy_0 (.O (d[0]), .CI (nx8473z1), .LI (nx8473z3)) ;
    XORCY xorcy_1 (.O (d[1]), .CI (nx8474z1), .LI (nx8474z2)) ;
    XORCY xorcy_2 (.O (d[2]), .CI (nx8475z1), .LI (nx8475z2)) ;
    XORCY xorcy_3 (.O (d[3]), .CI (nx8476z1), .LI (nx8476z2)) ;
    XORCY xorcy_4 (.O (d[4]), .CI (nx8477z1), .LI (nx8477z2)) ;
    XORCY xorcy_5 (.O (d[5]), .CI (nx8478z1), .LI (nx8478z2)) ;
    XORCY xorcy_6 (.O (d[6]), .CI (nx8479z1), .LI (nx8479z2)) ;
    XORCY xorcy_7 (.O (d[7]), .CI (nx8480z1), .LI (nx8480z2)) ;
    XORCY xorcy_8 (.O (d[8]), .CI (nx8481z1), .LI (nx8481z2)) ;
    XORCY xorcy_9 (.O (d[9]), .CI (nx8482z1), .LI (nx8482z2)) ;
    XORCY xorcy_10 (.O (d[10]), .CI (nx60018z1), .LI (nx60018z2)) ;
    XORCY xorcy_11 (.O (d[11]), .CI (nx60019z1), .LI (nx60019z2)) ;
    XORCY xorcy_12 (.O (d[12]), .CI (nx60020z1), .LI (nx60020z2)) ;
    XORCY xorcy_13 (.O (d[13]), .CI (nx60021z1), .LI (nx60021z2)) ;
    XORCY xorcy_14 (.O (d[14]), .CI (nx60022z1), .LI (nx60022z2)) ;
    XORCY xorcy_15 (.O (d[15]), .CI (nx60023z1), .LI (nx60023z2)) ;
    XORCY xorcy_16 (.O (d[16]), .CI (nx60024z1), .LI (nx60024z2)) ;
    XORCY xorcy_17 (.O (d[17]), .CI (nx60025z1), .LI (nx60025z2)) ;
    XORCY xorcy_18 (.O (d[18]), .CI (nx60026z1), .LI (nx60026z2)) ;
    XORCY xorcy_19 (.O (d[19]), .CI (nx60027z1), .LI (nx60027z2)) ;
    XORCY xorcy_20 (.O (d[20]), .CI (nx61015z1), .LI (nx61015z2)) ;
    XORCY xorcy_21 (.O (d[21]), .CI (nx61016z1), .LI (nx61016z2)) ;
    XORCY xorcy_22 (.O (d[22]), .CI (nx61017z1), .LI (nx61017z2)) ;
    XORCY xorcy_23 (.O (d[23]), .CI (nx61018z1), .LI (nx61018z2)) ;
    XORCY xorcy_24 (.O (d[24]), .CI (nx61019z1), .LI (nx61019z2)) ;
    XORCY xorcy_25 (.O (d[25]), .CI (nx61020z1), .LI (nx61020z2)) ;
    XORCY xorcy_26 (.O (d[26]), .CI (nx61021z1), .LI (nx61021z2)) ;
    XORCY xorcy_27 (.O (d[27]), .CI (nx61022z1), .LI (nx61022z2)) ;
    XORCY xorcy_28 (.O (d[28]), .CI (nx61023z1), .LI (nx61023z2)) ;
    XORCY xorcy_29 (.O (d[29]), .CI (nx19589z1), .LI (a[29])) ;
    LUT1 ix8473z1318 (.O (nx8473z3), .I0 (a[0])) ;
         defparam ix8473z1318.INIT = 4'h2;
    LUT1 ix8474z1316 (.O (nx8474z2), .I0 (a[1])) ;
         defparam ix8474z1316.INIT = 4'h2;
    LUT1 ix8475z1316 (.O (nx8475z2), .I0 (a[2])) ;
         defparam ix8475z1316.INIT = 4'h2;
    LUT1 ix8476z1316 (.O (nx8476z2), .I0 (a[3])) ;
         defparam ix8476z1316.INIT = 4'h2;
    LUT1 ix8477z1316 (.O (nx8477z2), .I0 (a[4])) ;
         defparam ix8477z1316.INIT = 4'h2;
    LUT1 ix8478z1316 (.O (nx8478z2), .I0 (a[5])) ;
         defparam ix8478z1316.INIT = 4'h2;
    LUT1 ix8479z1316 (.O (nx8479z2), .I0 (a[6])) ;
         defparam ix8479z1316.INIT = 4'h2;
    LUT1 ix8480z1316 (.O (nx8480z2), .I0 (a[7])) ;
         defparam ix8480z1316.INIT = 4'h2;
    LUT1 ix8481z1316 (.O (nx8481z2), .I0 (a[8])) ;
         defparam ix8481z1316.INIT = 4'h2;
    LUT1 ix8482z1316 (.O (nx8482z2), .I0 (a[9])) ;
         defparam ix8482z1316.INIT = 4'h2;
    LUT1 ix60018z1316 (.O (nx60018z2), .I0 (a[10])) ;
         defparam ix60018z1316.INIT = 4'h2;
    LUT1 ix60019z1316 (.O (nx60019z2), .I0 (a[11])) ;
         defparam ix60019z1316.INIT = 4'h2;
    LUT1 ix60020z1316 (.O (nx60020z2), .I0 (a[12])) ;
         defparam ix60020z1316.INIT = 4'h2;
    LUT1 ix60021z1316 (.O (nx60021z2), .I0 (a[13])) ;
         defparam ix60021z1316.INIT = 4'h2;
    LUT1 ix60022z1316 (.O (nx60022z2), .I0 (a[14])) ;
         defparam ix60022z1316.INIT = 4'h2;
    LUT1 ix60023z1316 (.O (nx60023z2), .I0 (a[15])) ;
         defparam ix60023z1316.INIT = 4'h2;
    LUT1 ix60024z1316 (.O (nx60024z2), .I0 (a[16])) ;
         defparam ix60024z1316.INIT = 4'h2;
    LUT1 ix60025z1316 (.O (nx60025z2), .I0 (a[17])) ;
         defparam ix60025z1316.INIT = 4'h2;
    LUT1 ix60026z1316 (.O (nx60026z2), .I0 (a[18])) ;
         defparam ix60026z1316.INIT = 4'h2;
    LUT1 ix60027z1316 (.O (nx60027z2), .I0 (a[19])) ;
         defparam ix60027z1316.INIT = 4'h2;
    LUT1 ix61015z1316 (.O (nx61015z2), .I0 (a[20])) ;
         defparam ix61015z1316.INIT = 4'h2;
    LUT1 ix61016z1316 (.O (nx61016z2), .I0 (a[21])) ;
         defparam ix61016z1316.INIT = 4'h2;
    LUT1 ix61017z1316 (.O (nx61017z2), .I0 (a[22])) ;
         defparam ix61017z1316.INIT = 4'h2;
    LUT1 ix61018z1316 (.O (nx61018z2), .I0 (a[23])) ;
         defparam ix61018z1316.INIT = 4'h2;
    LUT1 ix61019z1316 (.O (nx61019z2), .I0 (a[24])) ;
         defparam ix61019z1316.INIT = 4'h2;
    LUT1 ix61020z1316 (.O (nx61020z2), .I0 (a[25])) ;
         defparam ix61020z1316.INIT = 4'h2;
    LUT1 ix61021z1316 (.O (nx61021z2), .I0 (a[26])) ;
         defparam ix61021z1316.INIT = 4'h2;
    LUT1 ix61022z1316 (.O (nx61022z2), .I0 (a[27])) ;
         defparam ix61022z1316.INIT = 4'h2;
    LUT1 ix61023z1316 (.O (nx61023z2), .I0 (a[28])) ;
         defparam ix61023z1316.INIT = 4'h2;
    MUXCY muxcy_0 (.O (nx8474z1), .CI (nx8473z1), .DI (nx8473z2), .S (nx8473z3)
          ) ;
    MUXCY muxcy_1 (.O (nx8475z1), .CI (nx8474z1), .DI (nx8473z2), .S (nx8474z2)
          ) ;
    MUXCY muxcy_2 (.O (nx8476z1), .CI (nx8475z1), .DI (nx8473z2), .S (nx8475z2)
          ) ;
    MUXCY muxcy_3 (.O (nx8477z1), .CI (nx8476z1), .DI (nx8473z2), .S (nx8476z2)
          ) ;
    MUXCY muxcy_4 (.O (nx8478z1), .CI (nx8477z1), .DI (nx8473z2), .S (nx8477z2)
          ) ;
    MUXCY muxcy_5 (.O (nx8479z1), .CI (nx8478z1), .DI (nx8473z2), .S (nx8478z2)
          ) ;
    MUXCY muxcy_6 (.O (nx8480z1), .CI (nx8479z1), .DI (nx8473z2), .S (nx8479z2)
          ) ;
    MUXCY muxcy_7 (.O (nx8481z1), .CI (nx8480z1), .DI (nx8473z2), .S (nx8480z2)
          ) ;
    MUXCY muxcy_8 (.O (nx8482z1), .CI (nx8481z1), .DI (nx8473z2), .S (nx8481z2)
          ) ;
    MUXCY muxcy_9 (.O (nx60018z1), .CI (nx8482z1), .DI (nx8473z2), .S (nx8482z2)
          ) ;
    MUXCY muxcy_10 (.O (nx60019z1), .CI (nx60018z1), .DI (nx8473z2), .S (
          nx60018z2)) ;
    MUXCY muxcy_11 (.O (nx60020z1), .CI (nx60019z1), .DI (nx8473z2), .S (
          nx60019z2)) ;
    MUXCY muxcy_12 (.O (nx60021z1), .CI (nx60020z1), .DI (nx8473z2), .S (
          nx60020z2)) ;
    MUXCY muxcy_13 (.O (nx60022z1), .CI (nx60021z1), .DI (nx8473z2), .S (
          nx60021z2)) ;
    MUXCY muxcy_14 (.O (nx60023z1), .CI (nx60022z1), .DI (nx8473z2), .S (
          nx60022z2)) ;
    MUXCY muxcy_15 (.O (nx60024z1), .CI (nx60023z1), .DI (nx8473z2), .S (
          nx60023z2)) ;
    MUXCY muxcy_16 (.O (nx60025z1), .CI (nx60024z1), .DI (nx8473z2), .S (
          nx60024z2)) ;
    MUXCY muxcy_17 (.O (nx60026z1), .CI (nx60025z1), .DI (nx8473z2), .S (
          nx60025z2)) ;
    MUXCY muxcy_18 (.O (nx60027z1), .CI (nx60026z1), .DI (nx8473z2), .S (
          nx60026z2)) ;
    MUXCY muxcy_19 (.O (nx61015z1), .CI (nx60027z1), .DI (nx8473z2), .S (
          nx60027z2)) ;
    MUXCY muxcy_20 (.O (nx61016z1), .CI (nx61015z1), .DI (nx8473z2), .S (
          nx61015z2)) ;
    MUXCY muxcy_21 (.O (nx61017z1), .CI (nx61016z1), .DI (nx8473z2), .S (
          nx61016z2)) ;
    MUXCY muxcy_22 (.O (nx61018z1), .CI (nx61017z1), .DI (nx8473z2), .S (
          nx61017z2)) ;
    MUXCY muxcy_23 (.O (nx61019z1), .CI (nx61018z1), .DI (nx8473z2), .S (
          nx61018z2)) ;
    MUXCY muxcy_24 (.O (nx61020z1), .CI (nx61019z1), .DI (nx8473z2), .S (
          nx61019z2)) ;
    MUXCY muxcy_25 (.O (nx61021z1), .CI (nx61020z1), .DI (nx8473z2), .S (
          nx61020z2)) ;
    MUXCY muxcy_26 (.O (nx61022z1), .CI (nx61021z1), .DI (nx8473z2), .S (
          nx61021z2)) ;
    MUXCY muxcy_27 (.O (nx61023z1), .CI (nx61022z1), .DI (nx8473z2), .S (
          nx61022z2)) ;
    MUXCY muxcy_28 (.O (nx19589z1), .CI (nx61023z1), .DI (nx8473z2), .S (
          nx61023z2)) ;
endmodule


module ram_dq_32_1 ( wr_data1, rd_data1, addr1, wr_clk1, rd_clk1, wr_ena1, 
                     rd_ena1, ena1, rst1, regce1, regrst1, rd_access1, wr_data2, 
                     rd_data2, addr2, wr_clk2, rd_clk2, wr_ena2, rd_ena2, ena2, 
                     rst2, regce2, regrst2, rd_access2 ) ;

    input [31:0]wr_data1 ;
    output [31:0]rd_data1 ;
    input [4:0]addr1 ;
    input wr_clk1 ;
    input rd_clk1 ;
    input wr_ena1 ;
    input rd_ena1 ;
    input ena1 ;
    input rst1 ;
    input regce1 ;
    input regrst1 ;
    output rd_access1 ;
    input [31:0]wr_data2 ;
    output [31:0]rd_data2 ;
    input [4:0]addr2 ;
    input wr_clk2 ;
    input rd_clk2 ;
    input wr_ena2 ;
    input rd_ena2 ;
    input ena2 ;
    input rst2 ;
    input regce2 ;
    input regrst2 ;
    output rd_access2 ;




    RAM32M ROM_1 (.DOA ({rd_data2[1],rd_data2[0]}), .DOB ({rd_data2[3],
           rd_data2[2]}), .DOC ({rd_data2[5],rd_data2[4]}), .DOD ({rd_data2[7],
           rd_data2[6]}), .ADDRA ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}
           ), .ADDRB ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), .ADDRC ({
           addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), .ADDRD ({addr1[4],
           addr1[3],addr1[2],addr1[1],addr1[0]}), .DIA ({wr_data1[1],wr_data1[0]
           }), .DIB ({wr_data1[3],wr_data1[2]}), .DIC ({wr_data1[5],wr_data1[4]}
           ), .DID ({wr_data1[7],wr_data1[6]}), .WCLK (wr_clk1), .WE (wr_ena1)
           ) ;
    RAM32M ROM_2 (.DOA ({rd_data2[9],rd_data2[8]}), .DOB ({rd_data2[11],
           rd_data2[10]}), .DOC ({rd_data2[13],rd_data2[12]}), .DOD ({
           rd_data2[15],rd_data2[14]}), .ADDRA ({addr1[4],addr1[3],addr1[2],
           addr1[1],addr1[0]}), .ADDRB ({addr1[4],addr1[3],addr1[2],addr1[1],
           addr1[0]}), .ADDRC ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), 
           .ADDRD ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), .DIA ({
           wr_data1[9],wr_data1[8]}), .DIB ({wr_data1[11],wr_data1[10]}), .DIC (
           {wr_data1[13],wr_data1[12]}), .DID ({wr_data1[15],wr_data1[14]}), .WCLK (
           wr_clk1), .WE (wr_ena1)) ;
    RAM32M ROM_3 (.DOA ({rd_data2[17],rd_data2[16]}), .DOB ({rd_data2[19],
           rd_data2[18]}), .DOC ({rd_data2[21],rd_data2[20]}), .DOD ({
           rd_data2[23],rd_data2[22]}), .ADDRA ({addr1[4],addr1[3],addr1[2],
           addr1[1],addr1[0]}), .ADDRB ({addr1[4],addr1[3],addr1[2],addr1[1],
           addr1[0]}), .ADDRC ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), 
           .ADDRD ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), .DIA ({
           wr_data1[17],wr_data1[16]}), .DIB ({wr_data1[19],wr_data1[18]}), .DIC (
           {wr_data1[21],wr_data1[20]}), .DID ({wr_data1[23],wr_data1[22]}), .WCLK (
           wr_clk1), .WE (wr_ena1)) ;
    RAM32M ROM_4 (.DOA ({rd_data2[25],rd_data2[24]}), .DOB ({rd_data2[27],
           rd_data2[26]}), .DOC ({rd_data2[29],rd_data2[28]}), .DOD ({
           rd_data2[31],rd_data2[30]}), .ADDRA ({addr1[4],addr1[3],addr1[2],
           addr1[1],addr1[0]}), .ADDRB ({addr1[4],addr1[3],addr1[2],addr1[1],
           addr1[0]}), .ADDRC ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), 
           .ADDRD ({addr1[4],addr1[3],addr1[2],addr1[1],addr1[0]}), .DIA ({
           wr_data1[25],wr_data1[24]}), .DIB ({wr_data1[27],wr_data1[26]}), .DIC (
           {wr_data1[29],wr_data1[28]}), .DID ({wr_data1[31],wr_data1[30]}), .WCLK (
           wr_clk1), .WE (wr_ena1)) ;
endmodule


module ram_dq_32_0 ( wr_data1, rd_data1, addr1, wr_clk1, rd_clk1, wr_ena1, 
                     rd_ena1, ena1, rst1, regce1, regrst1, rd_access1, wr_data2, 
                     rd_data2, addr2, wr_clk2, rd_clk2, wr_ena2, rd_ena2, ena2, 
                     rst2, regce2, regrst2, rd_access2, wr_data3, rd_data3, 
                     addr3, wr_clk3, rd_clk3, wr_ena3, rd_ena3, ena3, rst3, 
                     regce3, regrst3, rd_access3 ) ;

    input [31:0]wr_data1 ;
    output [31:0]rd_data1 ;
    input [4:0]addr1 ;
    input wr_clk1 ;
    input rd_clk1 ;
    input wr_ena1 ;
    input rd_ena1 ;
    input ena1 ;
    input rst1 ;
    input regce1 ;
    input regrst1 ;
    output rd_access1 ;
    input [31:0]wr_data2 ;
    output [31:0]rd_data2 ;
    input [4:0]addr2 ;
    input wr_clk2 ;
    input rd_clk2 ;
    input wr_ena2 ;
    input rd_ena2 ;
    input ena2 ;
    input rst2 ;
    input regce2 ;
    input regrst2 ;
    output rd_access2 ;
    input [31:0]wr_data3 ;
    output [31:0]rd_data3 ;
    input [4:0]addr3 ;
    input wr_clk3 ;
    input rd_clk3 ;
    input wr_ena3 ;
    input rd_ena3 ;
    input ena3 ;
    input rst3 ;
    input regce3 ;
    input regrst3 ;
    output rd_access3 ;

    wire [3:0]addr1_rename3;
    wire [23:0] \$dummy ;




    GND ps_gnd (.G (addr1_rename3[3])) ;
    RAM32M register_1 (.DOA ({rd_data2[1],rd_data2[0]}), .DOB ({rd_data2[3],
           rd_data2[2]}), .DOC ({rd_data2[5],rd_data2[4]}), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[1],wr_data1[0]}), .DIB ({wr_data1[3],wr_data1[2]}), .DIC ({
           wr_data1[5],wr_data1[4]}), .DID ({addr1_rename3[3],addr1_rename3[3]})
           , .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_2 (.DOA ({rd_data2[7],rd_data2[6]}), .DOB ({rd_data2[9],
           rd_data2[8]}), .DOC ({rd_data2[11],rd_data2[10]}), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[7],wr_data1[6]}), .DIB ({wr_data1[9],wr_data1[8]}), .DIC ({
           wr_data1[11],wr_data1[10]}), .DID ({addr1_rename3[3],addr1_rename3[3]
           }), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_3 (.DOA ({rd_data2[13],rd_data2[12]}), .DOB ({rd_data2[15],
           rd_data2[14]}), .DOC ({rd_data2[17],rd_data2[16]}), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[13],wr_data1[12]}), .DIB ({wr_data1[15],wr_data1[14]}), .DIC (
           {wr_data1[17],wr_data1[16]}), .DID ({addr1_rename3[3],
           addr1_rename3[3]}), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_4 (.DOA ({rd_data2[19],rd_data2[18]}), .DOB ({rd_data2[21],
           rd_data2[20]}), .DOC ({rd_data2[23],rd_data2[22]}), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[19],wr_data1[18]}), .DIB ({wr_data1[21],wr_data1[20]}), .DIC (
           {wr_data1[23],wr_data1[22]}), .DID ({addr1_rename3[3],
           addr1_rename3[3]}), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_5 (.DOA ({rd_data2[25],rd_data2[24]}), .DOB ({rd_data2[27],
           rd_data2[26]}), .DOC ({rd_data2[29],rd_data2[28]}), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[25],wr_data1[24]}), .DIB ({wr_data1[27],wr_data1[26]}), .DIC (
           {wr_data1[29],wr_data1[28]}), .DID ({addr1_rename3[3],
           addr1_rename3[3]}), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM64M register_6 (.DOA (rd_data2[30]), .DOB (rd_data2[31]), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],
           addr2[0]}), .ADDRB ({addr1_rename3[3],addr1_rename3[3],
           addr1_rename3[3],addr2[2],addr2[1],addr2[0]}), .ADDRC ({
           addr1_rename3[3],addr1_rename3[3],addr1_rename3[3],addr2[2],addr2[1],
           addr2[0]}), .ADDRD ({addr1_rename3[3],addr1_rename3[3],
           addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (wr_data1[30]), .DIB (
           wr_data1[31]), .DIC (addr1_rename3[3]), .DID (addr1_rename3[3]), .WCLK (
           wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_1_1_0 (.DOA ({rd_data3[1],rd_data3[0]}), .DOB ({rd_data3[3],
           rd_data3[2]}), .DOC ({rd_data3[5],rd_data3[4]}), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[1],wr_data1[0]}), .DIB ({wr_data1[3],wr_data1[2]}), .DIC ({
           wr_data1[5],wr_data1[4]}), .DID ({addr1_rename3[3],addr1_rename3[3]})
           , .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_2_1_0 (.DOA ({rd_data3[7],rd_data3[6]}), .DOB ({rd_data3[9],
           rd_data3[8]}), .DOC ({rd_data3[11],rd_data3[10]}), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[7],wr_data1[6]}), .DIB ({wr_data1[9],wr_data1[8]}), .DIC ({
           wr_data1[11],wr_data1[10]}), .DID ({addr1_rename3[3],addr1_rename3[3]
           }), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_3_1_0 (.DOA ({rd_data3[13],rd_data3[12]}), .DOB ({
           rd_data3[15],rd_data3[14]}), .DOC ({rd_data3[17],rd_data3[16]}), .ADDRA (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[13],wr_data1[12]}), .DIB ({wr_data1[15],wr_data1[14]}), .DIC (
           {wr_data1[17],wr_data1[16]}), .DID ({addr1_rename3[3],
           addr1_rename3[3]}), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_4_1_0 (.DOA ({rd_data3[19],rd_data3[18]}), .DOB ({
           rd_data3[21],rd_data3[20]}), .DOC ({rd_data3[23],rd_data3[22]}), .ADDRA (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[19],wr_data1[18]}), .DIB ({wr_data1[21],wr_data1[20]}), .DIC (
           {wr_data1[23],wr_data1[22]}), .DID ({addr1_rename3[3],
           addr1_rename3[3]}), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM32M register_5_1_0 (.DOA ({rd_data3[25],rd_data3[24]}), .DOB ({
           rd_data3[27],rd_data3[26]}), .DOC ({rd_data3[29],rd_data3[28]}), .ADDRA (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRB (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRC (
           {addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRD (
           {addr1_rename3[3],addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (
           {wr_data1[25],wr_data1[24]}), .DIB ({wr_data1[27],wr_data1[26]}), .DIC (
           {wr_data1[29],wr_data1[28]}), .DID ({addr1_rename3[3],
           addr1_rename3[3]}), .WCLK (wr_clk1), .WE (wr_ena1)) ;
    RAM64M register_6_1_0 (.DOA (rd_data3[30]), .DOB (rd_data3[31]), .ADDRA ({
           addr1_rename3[3],addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],
           addr3[0]}), .ADDRB ({addr1_rename3[3],addr1_rename3[3],
           addr1_rename3[3],addr3[2],addr3[1],addr3[0]}), .ADDRC ({
           addr1_rename3[3],addr1_rename3[3],addr1_rename3[3],addr3[2],addr3[1],
           addr3[0]}), .ADDRD ({addr1_rename3[3],addr1_rename3[3],
           addr1_rename3[3],addr1[2],addr1[1],addr1[0]}), .DIA (wr_data1[30]), .DIB (
           wr_data1[31]), .DIC (addr1_rename3[3]), .DID (addr1_rename3[3]), .WCLK (
           wr_clk1), .WE (wr_ena1)) ;
endmodule

